// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition"

// DATE "06/11/2023 10:37:46"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module IFFT (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk,
	reset_n,
	sink_valid,
	sink_ready,
	sink_error,
	sink_sop,
	sink_eop,
	sink_real,
	sink_imag,
	inverse,
	source_valid,
	source_ready,
	source_error,
	source_sop,
	source_eop,
	source_real,
	source_imag,
	source_exp)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk;
input 	reset_n;
input 	sink_valid;
output 	sink_ready;
input 	[1:0] sink_error;
input 	sink_sop;
input 	sink_eop;
input 	[7:0] sink_real;
input 	[7:0] sink_imag;
input 	[0:0] inverse;
output 	source_valid;
input 	source_ready;
output 	[1:0] source_error;
output 	source_sop;
output 	source_eop;
output 	[7:0] source_real;
output 	[7:0] source_imag;
output 	[5:0] source_exp;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;
wire \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;
wire \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;
wire \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;
wire \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;
wire \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;
wire \fft_ii_0|source_real[0]~combout ;
wire \fft_ii_0|source_real[1]~combout ;
wire \fft_ii_0|source_real[2]~combout ;
wire \fft_ii_0|source_real[3]~combout ;
wire \fft_ii_0|source_real[4]~combout ;
wire \fft_ii_0|source_real[5]~combout ;
wire \fft_ii_0|source_real[6]~combout ;
wire \fft_ii_0|source_real[7]~combout ;
wire \fft_ii_0|source_imag[0]~combout ;
wire \fft_ii_0|source_imag[1]~combout ;
wire \fft_ii_0|source_imag[2]~combout ;
wire \fft_ii_0|source_imag[3]~combout ;
wire \fft_ii_0|source_imag[4]~combout ;
wire \fft_ii_0|source_imag[5]~combout ;
wire \fft_ii_0|source_imag[6]~combout ;
wire \fft_ii_0|source_imag[7]~combout ;
wire \fft_ii_0|source_exp[0]~combout ;
wire \fft_ii_0|source_exp[1]~combout ;
wire \fft_ii_0|source_exp[2]~combout ;
wire \fft_ii_0|source_exp[3]~combout ;
wire \fft_ii_0|source_exp[4]~combout ;
wire \fft_ii_0|source_exp[5]~combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \source_ready~input_o ;
wire \sink_eop~input_o ;
wire \sink_valid~input_o ;
wire \sink_error[0]~input_o ;
wire \sink_error[1]~input_o ;
wire \sink_sop~input_o ;
wire \inverse[0]~input_o ;
wire \sink_real[6]~input_o ;
wire \sink_imag[6]~input_o ;
wire \sink_real[5]~input_o ;
wire \sink_imag[5]~input_o ;
wire \sink_real[2]~input_o ;
wire \sink_imag[2]~input_o ;
wire \sink_real[3]~input_o ;
wire \sink_imag[3]~input_o ;
wire \sink_real[4]~input_o ;
wire \sink_imag[4]~input_o ;
wire \sink_real[7]~input_o ;
wire \sink_imag[7]~input_o ;
wire \sink_real[0]~input_o ;
wire \sink_imag[0]~input_o ;
wire \sink_real[1]~input_o ;
wire \sink_imag[1]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ;
wire \nabboc|pzdyqx_impl_inst|sdr~combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


IFFT_IFFT_fft_ii_0 fft_ii_0(
	.at_sink_ready_s(\fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ),
	.at_source_valid_s(\fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ),
	.at_source_error_0(\fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ),
	.at_source_error_1(\fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ),
	.at_source_sop_s(\fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ),
	.at_source_eop_s(\fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ),
	.source_real_0(\fft_ii_0|source_real[0]~combout ),
	.source_real_1(\fft_ii_0|source_real[1]~combout ),
	.source_real_2(\fft_ii_0|source_real[2]~combout ),
	.source_real_3(\fft_ii_0|source_real[3]~combout ),
	.source_real_4(\fft_ii_0|source_real[4]~combout ),
	.source_real_5(\fft_ii_0|source_real[5]~combout ),
	.source_real_6(\fft_ii_0|source_real[6]~combout ),
	.source_real_7(\fft_ii_0|source_real[7]~combout ),
	.source_imag_0(\fft_ii_0|source_imag[0]~combout ),
	.source_imag_1(\fft_ii_0|source_imag[1]~combout ),
	.source_imag_2(\fft_ii_0|source_imag[2]~combout ),
	.source_imag_3(\fft_ii_0|source_imag[3]~combout ),
	.source_imag_4(\fft_ii_0|source_imag[4]~combout ),
	.source_imag_5(\fft_ii_0|source_imag[5]~combout ),
	.source_imag_6(\fft_ii_0|source_imag[6]~combout ),
	.source_imag_7(\fft_ii_0|source_imag[7]~combout ),
	.source_exp_0(\fft_ii_0|source_exp[0]~combout ),
	.source_exp_1(\fft_ii_0|source_exp[1]~combout ),
	.source_exp_2(\fft_ii_0|source_exp[2]~combout ),
	.source_exp_3(\fft_ii_0|source_exp[3]~combout ),
	.source_exp_4(\fft_ii_0|source_exp[4]~combout ),
	.source_exp_5(\fft_ii_0|source_exp[5]~combout ),
	.GND_port(\~GND~combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.source_ready(\source_ready~input_o ),
	.sink_eop(\sink_eop~input_o ),
	.sink_valid(\sink_valid~input_o ),
	.sink_error_0(\sink_error[0]~input_o ),
	.sink_error_1(\sink_error[1]~input_o ),
	.sink_sop(\sink_sop~input_o ),
	.inverse_0(\inverse[0]~input_o ),
	.sink_real_6(\sink_real[6]~input_o ),
	.sink_imag_6(\sink_imag[6]~input_o ),
	.sink_real_5(\sink_real[5]~input_o ),
	.sink_imag_5(\sink_imag[5]~input_o ),
	.sink_real_2(\sink_real[2]~input_o ),
	.sink_imag_2(\sink_imag[2]~input_o ),
	.sink_real_3(\sink_real[3]~input_o ),
	.sink_imag_3(\sink_imag[3]~input_o ),
	.sink_real_4(\sink_real[4]~input_o ),
	.sink_imag_4(\sink_imag[4]~input_o ),
	.sink_real_7(\sink_real[7]~input_o ),
	.sink_imag_7(\sink_imag[7]~input_o ),
	.sink_real_0(\sink_real[0]~input_o ),
	.sink_imag_0(\sink_imag[0]~input_o ),
	.sink_real_1(\sink_real[1]~input_o ),
	.sink_imag_1(\sink_imag[1]~input_o ));

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \source_ready~input_o  = source_ready;

assign \sink_eop~input_o  = sink_eop;

assign \sink_valid~input_o  = sink_valid;

assign \sink_error[0]~input_o  = sink_error[0];

assign \sink_error[1]~input_o  = sink_error[1];

assign \sink_sop~input_o  = sink_sop;

assign \inverse[0]~input_o  = inverse[0];

assign \sink_real[6]~input_o  = sink_real[6];

assign \sink_imag[6]~input_o  = sink_imag[6];

assign \sink_real[5]~input_o  = sink_real[5];

assign \sink_imag[5]~input_o  = sink_imag[5];

assign \sink_real[2]~input_o  = sink_real[2];

assign \sink_imag[2]~input_o  = sink_imag[2];

assign \sink_real[3]~input_o  = sink_real[3];

assign \sink_imag[3]~input_o  = sink_imag[3];

assign \sink_real[4]~input_o  = sink_real[4];

assign \sink_imag[4]~input_o  = sink_imag[4];

assign \sink_real[7]~input_o  = sink_real[7];

assign \sink_imag[7]~input_o  = sink_imag[7];

assign \sink_real[0]~input_o  = sink_real[0];

assign \sink_imag[0]~input_o  = sink_imag[0];

assign \sink_real[1]~input_o  = sink_real[1];

assign \sink_imag[1]~input_o  = sink_imag[1];

assign sink_ready = \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_sink_1|at_sink_ready_s~q ;

assign source_valid = \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_valid_s~q ;

assign source_error[0] = \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_error[0]~q ;

assign source_error[1] = \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_error[1]~q ;

assign source_sop = \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_sop_s~q ;

assign source_eop = \fft_ii_0|asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_eop_s~q ;

assign source_real[0] = \fft_ii_0|source_real[0]~combout ;

assign source_real[1] = \fft_ii_0|source_real[1]~combout ;

assign source_real[2] = \fft_ii_0|source_real[2]~combout ;

assign source_real[3] = \fft_ii_0|source_real[3]~combout ;

assign source_real[4] = \fft_ii_0|source_real[4]~combout ;

assign source_real[5] = \fft_ii_0|source_real[5]~combout ;

assign source_real[6] = \fft_ii_0|source_real[6]~combout ;

assign source_real[7] = \fft_ii_0|source_real[7]~combout ;

assign source_imag[0] = \fft_ii_0|source_imag[0]~combout ;

assign source_imag[1] = \fft_ii_0|source_imag[1]~combout ;

assign source_imag[2] = \fft_ii_0|source_imag[2]~combout ;

assign source_imag[3] = \fft_ii_0|source_imag[3]~combout ;

assign source_imag[4] = \fft_ii_0|source_imag[4]~combout ;

assign source_imag[5] = \fft_ii_0|source_imag[5]~combout ;

assign source_imag[6] = \fft_ii_0|source_imag[6]~combout ;

assign source_imag[7] = \fft_ii_0|source_imag[7]~combout ;

assign source_exp[0] = \fft_ii_0|source_exp[0]~combout ;

assign source_exp[1] = \fft_ii_0|source_exp[1]~combout ;

assign source_exp[2] = \fft_ii_0|source_exp[2]~combout ;

assign source_exp[3] = \fft_ii_0|source_exp[3]~combout ;

assign source_exp[4] = \fft_ii_0|source_exp[4]~combout ;

assign source_exp[5] = \fft_ii_0|source_exp[5]~combout ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\~GND~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFBF7FFFFF7FBFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'h7FFFDFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .lut_mask = 64'hDEDEDEDEDEDEDEDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .lut_mask = 64'hEDDEDEEDDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_1 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_2 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'hDFD5FFFFDFD5FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|AMGP4450~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|AMGP4450 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .lut_mask = 64'hBFFBFFFFBFFBFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .lut_mask = 64'hFF96FFF6FF96FFF6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .lut_mask = 64'hF9F6F9F6F9F6F9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .lut_mask = 64'h9F6FF9F69F6FF9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\altera_internal_jtag~TDIUTAP ),
	.dataf(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|sdr (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|sdr .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|sdr .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \nabboc|pzdyqx_impl_inst|sdr .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'hF0F0F0F0FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h0FF00FF0FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'hF00F0FF0FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'h5AA5A55AFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'h96696996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~4_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFAFFFAFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h5F3FFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hAFFAAFFAAFFAAFFA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hBEEBBEEBEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'hD8FFFFFFD8FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hEFFFFEFFEFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'hFF96FFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hF7FFFFFF37FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module IFFT_IFFT_fft_ii_0 (
	at_sink_ready_s,
	at_source_valid_s,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s,
	at_source_eop_s,
	source_real_0,
	source_real_1,
	source_real_2,
	source_real_3,
	source_real_4,
	source_real_5,
	source_real_6,
	source_real_7,
	source_imag_0,
	source_imag_1,
	source_imag_2,
	source_imag_3,
	source_imag_4,
	source_imag_5,
	source_imag_6,
	source_imag_7,
	source_exp_0,
	source_exp_1,
	source_exp_2,
	source_exp_3,
	source_exp_4,
	source_exp_5,
	GND_port,
	NJQG9082,
	clk,
	reset_n,
	source_ready,
	sink_eop,
	sink_valid,
	sink_error_0,
	sink_error_1,
	sink_sop,
	inverse_0,
	sink_real_6,
	sink_imag_6,
	sink_real_5,
	sink_imag_5,
	sink_real_2,
	sink_imag_2,
	sink_real_3,
	sink_imag_3,
	sink_real_4,
	sink_imag_4,
	sink_real_7,
	sink_imag_7,
	sink_real_0,
	sink_imag_0,
	sink_real_1,
	sink_imag_1)/* synthesis synthesis_greybox=1 */;
output 	at_sink_ready_s;
output 	at_source_valid_s;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s;
output 	at_source_eop_s;
output 	source_real_0;
output 	source_real_1;
output 	source_real_2;
output 	source_real_3;
output 	source_real_4;
output 	source_real_5;
output 	source_real_6;
output 	source_real_7;
output 	source_imag_0;
output 	source_imag_1;
output 	source_imag_2;
output 	source_imag_3;
output 	source_imag_4;
output 	source_imag_5;
output 	source_imag_6;
output 	source_imag_7;
output 	source_exp_0;
output 	source_exp_1;
output 	source_exp_2;
output 	source_exp_3;
output 	source_exp_4;
output 	source_exp_5;
input 	GND_port;
input 	NJQG9082;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_eop;
input 	sink_valid;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_sop;
input 	inverse_0;
input 	sink_real_6;
input 	sink_imag_6;
input 	sink_real_5;
input 	sink_imag_5;
input 	sink_real_2;
input 	sink_imag_2;
input 	sink_real_3;
input 	sink_imag_3;
input 	sink_real_4;
input 	sink_imag_4;
input 	sink_real_7;
input 	sink_imag_7;
input 	sink_real_0;
input 	sink_imag_0;
input 	sink_real_1;
input 	sink_imag_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ;
wire \asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ;


IFFT_asj_fft_sglstream asj_fft_sglstream_inst(
	.at_source_data_14(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ),
	.at_source_data_15(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ),
	.at_source_data_16(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ),
	.at_source_data_17(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ),
	.at_source_data_18(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ),
	.at_source_data_19(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ),
	.at_source_data_20(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ),
	.at_source_data_21(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ),
	.at_source_data_6(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ),
	.at_source_data_7(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ),
	.at_source_data_8(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ),
	.at_source_data_9(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ),
	.at_source_data_10(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ),
	.at_source_data_11(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ),
	.at_source_data_12(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ),
	.at_source_data_13(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ),
	.at_source_data_0(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ),
	.at_source_data_1(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ),
	.at_source_data_2(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ),
	.at_source_data_3(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ),
	.at_source_data_4(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ),
	.at_source_data_5(\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ),
	.at_sink_ready_s(at_sink_ready_s),
	.at_source_valid_s(at_source_valid_s),
	.at_source_error_0(at_source_error_0),
	.at_source_error_1(at_source_error_1),
	.at_source_sop_s(at_source_sop_s),
	.at_source_eop_s(at_source_eop_s),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready),
	.sink_eop(sink_eop),
	.sink_valid(sink_valid),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.sink_sop(sink_sop),
	.inverse_0(inverse_0),
	.sink_real({sink_real_7,sink_real_6,sink_real_5,sink_real_4,sink_real_3,sink_real_2,sink_real_1,sink_real_0}),
	.sink_imag({sink_imag_7,sink_imag_6,sink_imag_5,sink_imag_4,sink_imag_3,sink_imag_2,sink_imag_1,sink_imag_0}));

cyclonev_lcell_comb \source_real[0] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[0] .extended_lut = "off";
defparam \source_real[0] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[0] .shared_arith = "off";

cyclonev_lcell_comb \source_real[1] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[1] .extended_lut = "off";
defparam \source_real[1] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[1] .shared_arith = "off";

cyclonev_lcell_comb \source_real[2] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[2] .extended_lut = "off";
defparam \source_real[2] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[2] .shared_arith = "off";

cyclonev_lcell_comb \source_real[3] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[3] .extended_lut = "off";
defparam \source_real[3] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[3] .shared_arith = "off";

cyclonev_lcell_comb \source_real[4] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[4] .extended_lut = "off";
defparam \source_real[4] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[4] .shared_arith = "off";

cyclonev_lcell_comb \source_real[5] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[5] .extended_lut = "off";
defparam \source_real[5] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[5] .shared_arith = "off";

cyclonev_lcell_comb \source_real[6] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[6] .extended_lut = "off";
defparam \source_real[6] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[6] .shared_arith = "off";

cyclonev_lcell_comb \source_real[7] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_real_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_real[7] .extended_lut = "off";
defparam \source_real[7] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_real[7] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[0] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[0] .extended_lut = "off";
defparam \source_imag[0] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[0] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[1] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[1] .extended_lut = "off";
defparam \source_imag[1] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[1] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[2] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[2] .extended_lut = "off";
defparam \source_imag[2] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[2] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[3] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[3] .extended_lut = "off";
defparam \source_imag[3] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[3] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[4] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[4] .extended_lut = "off";
defparam \source_imag[4] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[4] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[5] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[5] .extended_lut = "off";
defparam \source_imag[5] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[5] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[6] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[6] .extended_lut = "off";
defparam \source_imag[6] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[6] .shared_arith = "off";

cyclonev_lcell_comb \source_imag[7] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_imag_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_imag[7] .extended_lut = "off";
defparam \source_imag[7] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_imag[7] .shared_arith = "off";

cyclonev_lcell_comb \source_exp[0] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_exp_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_exp[0] .extended_lut = "off";
defparam \source_exp[0] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_exp[0] .shared_arith = "off";

cyclonev_lcell_comb \source_exp[1] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_exp_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_exp[1] .extended_lut = "off";
defparam \source_exp[1] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_exp[1] .shared_arith = "off";

cyclonev_lcell_comb \source_exp[2] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_exp_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_exp[2] .extended_lut = "off";
defparam \source_exp[2] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_exp[2] .shared_arith = "off";

cyclonev_lcell_comb \source_exp[3] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_exp_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_exp[3] .extended_lut = "off";
defparam \source_exp[3] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_exp[3] .shared_arith = "off";

cyclonev_lcell_comb \source_exp[4] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_exp_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_exp[4] .extended_lut = "off";
defparam \source_exp[4] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_exp[4] .shared_arith = "off";

cyclonev_lcell_comb \source_exp[5] (
	.dataa(!NJQG9082),
	.datab(!\asj_fft_sglstream_inst|auk_dsp_atlantic_source_1|at_source_data[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(source_exp_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_exp[5] .extended_lut = "off";
defparam \source_exp[5] .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \source_exp[5] .shared_arith = "off";

endmodule

module IFFT_asj_fft_sglstream (
	at_source_data_14,
	at_source_data_15,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	at_sink_ready_s,
	at_source_valid_s,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s,
	at_source_eop_s,
	GND_port,
	clk,
	reset_n,
	source_ready,
	sink_eop,
	sink_valid,
	sink_error_0,
	sink_error_1,
	sink_sop,
	inverse_0,
	sink_real,
	sink_imag)/* synthesis synthesis_greybox=1 */;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
output 	at_sink_ready_s;
output 	at_source_valid_s;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s;
output 	at_source_eop_s;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_eop;
input 	sink_valid;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_sop;
input 	inverse_0;
input 	[7:0] sink_real;
input 	[7:0] sink_imag;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_in_work~q ;
wire \master_source_ena~q ;
wire \fft_real_out[0]~q ;
wire \fft_real_out[1]~q ;
wire \fft_real_out[2]~q ;
wire \fft_real_out[3]~q ;
wire \fft_real_out[4]~q ;
wire \fft_real_out[5]~q ;
wire \fft_real_out[6]~q ;
wire \fft_real_out[7]~q ;
wire \fft_imag_out[0]~q ;
wire \fft_imag_out[1]~q ;
wire \fft_imag_out[2]~q ;
wire \fft_imag_out[3]~q ;
wire \fft_imag_out[4]~q ;
wire \fft_imag_out[5]~q ;
wire \fft_imag_out[6]~q ;
wire \fft_imag_out[7]~q ;
wire \oe~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[0]~q ;
wire \fft_dirn_stream~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[1]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[2]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[3]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[4]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[5]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[6]~q ;
wire \gen_radix_4_last_pass:lpp|data_real_o[7]~q ;
wire \fft_s2_cur.WAIT_FOR_LPP_INPUT~q ;
wire \sop_out~q ;
wire \fft_dirn_held_o2~q ;
wire \lpp_count_offset[5]~q ;
wire \lpp_count_offset[1]~q ;
wire \lpp_count_offset[2]~q ;
wire \lpp_count_offset[3]~q ;
wire \lpp_count_offset[4]~q ;
wire \delay_lpp_en|tdl_arr[5]~q ;
wire \fft_dirn_held_o~q ;
wire \gen_le256_mk:ctrl|blk_done_int~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ;
wire \lpp_count[0]~q ;
wire \lpp_count[1]~q ;
wire \lpp_count[2]~q ;
wire \lpp_count[3]~q ;
wire \lpp_count[4]~q ;
wire \lpp_count[5]~q ;
wire \writer|next_block~q ;
wire \fft_dirn_held~q ;
wire \gen_le256_mk:ctrl|p[0]~q ;
wire \Add2~1_sumout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add2~9_sumout ;
wire \Add2~10 ;
wire \Add2~13_sumout ;
wire \Add2~14 ;
wire \Add2~17_sumout ;
wire \Add2~18 ;
wire \Add2~21_sumout ;
wire \fft_dirn~q ;
wire \data_rdy_vec[4]~q ;
wire \gen_le256_mk:ctrl|next_pass_i~q ;
wire \data_rdy_vec[3]~q ;
wire \gen_dft_1:delay_blk_done|tdl_arr[11]~q ;
wire \data_rdy_vec[2]~q ;
wire \data_rdy_vec[1]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][3]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][7]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][7]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][3]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][4]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][4]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][5]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][5]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][6]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][6]~q ;
wire \data_rdy_vec[0]~q ;
wire \gen_dft_1:delay_blk_done2|tdl_arr[19]~q ;
wire \writer|data_rdy_int~q ;
wire \lpp_ram_data_out[3][10]~q ;
wire \lpp_ram_data_out[0][10]~q ;
wire \lpp_ram_data_out[1][10]~q ;
wire \lpp_ram_data_out[2][10]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ;
wire \lpp_ram_data_out[3][2]~q ;
wire \lpp_ram_data_out[0][2]~q ;
wire \lpp_ram_data_out[1][2]~q ;
wire \lpp_ram_data_out[2][2]~q ;
wire \lpp_ram_data_out[3][11]~q ;
wire \lpp_ram_data_out[0][11]~q ;
wire \lpp_ram_data_out[1][11]~q ;
wire \lpp_ram_data_out[2][11]~q ;
wire \lpp_ram_data_out[3][3]~q ;
wire \lpp_ram_data_out[0][3]~q ;
wire \lpp_ram_data_out[1][3]~q ;
wire \lpp_ram_data_out[2][3]~q ;
wire \lpp_ram_data_out[3][12]~q ;
wire \lpp_ram_data_out[0][12]~q ;
wire \lpp_ram_data_out[1][12]~q ;
wire \lpp_ram_data_out[2][12]~q ;
wire \lpp_ram_data_out[3][4]~q ;
wire \lpp_ram_data_out[0][4]~q ;
wire \lpp_ram_data_out[1][4]~q ;
wire \lpp_ram_data_out[2][4]~q ;
wire \lpp_ram_data_out[3][13]~q ;
wire \lpp_ram_data_out[0][13]~q ;
wire \lpp_ram_data_out[1][13]~q ;
wire \lpp_ram_data_out[2][13]~q ;
wire \lpp_ram_data_out[3][5]~q ;
wire \lpp_ram_data_out[0][5]~q ;
wire \lpp_ram_data_out[1][5]~q ;
wire \lpp_ram_data_out[2][5]~q ;
wire \lpp_ram_data_out[3][14]~q ;
wire \lpp_ram_data_out[0][14]~q ;
wire \lpp_ram_data_out[1][14]~q ;
wire \lpp_ram_data_out[2][14]~q ;
wire \lpp_ram_data_out[3][6]~q ;
wire \lpp_ram_data_out[0][6]~q ;
wire \lpp_ram_data_out[1][6]~q ;
wire \lpp_ram_data_out[2][6]~q ;
wire \lpp_ram_data_out[3][15]~q ;
wire \lpp_ram_data_out[0][15]~q ;
wire \lpp_ram_data_out[1][15]~q ;
wire \lpp_ram_data_out[2][15]~q ;
wire \lpp_ram_data_out[3][7]~q ;
wire \lpp_ram_data_out[0][7]~q ;
wire \lpp_ram_data_out[1][7]~q ;
wire \lpp_ram_data_out[2][7]~q ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \lpp_sel~q ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \lpp_ram_data_out[3][9]~q ;
wire \lpp_ram_data_out[0][9]~q ;
wire \lpp_ram_data_out[1][9]~q ;
wire \lpp_ram_data_out[2][9]~q ;
wire \lpp_ram_data_out[3][1]~q ;
wire \lpp_ram_data_out[0][1]~q ;
wire \lpp_ram_data_out[1][1]~q ;
wire \lpp_ram_data_out[2][1]~q ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \wc_vec[3]~q ;
wire \gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ;
wire \gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ;
wire \rdaddress_c_bus[0]~q ;
wire \rdaddress_c_bus[13]~q ;
wire \rdaddress_c_bus[10]~q ;
wire \rdaddress_c_bus[3]~q ;
wire \wd_vec[3]~q ;
wire \rdaddress_c_bus[14]~q ;
wire \rdaddress_c_bus[15]~q ;
wire \rdaddress_c_bus[11]~q ;
wire \rdaddress_c_bus[7]~q ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \lpp_ram_data_out[3][8]~q ;
wire \lpp_ram_data_out[0][8]~q ;
wire \lpp_ram_data_out[1][8]~q ;
wire \lpp_ram_data_out[2][8]~q ;
wire \lpp_ram_data_out[3][0]~q ;
wire \lpp_ram_data_out[0][0]~q ;
wire \lpp_ram_data_out[1][0]~q ;
wire \lpp_ram_data_out[2][0]~q ;
wire \wc_vec[2]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][2]~q ;
wire \gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a3~portbdataout ;
wire \gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a2~portbdataout ;
wire \gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ;
wire \gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ;
wire \wd_vec[2]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][2]~q ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \wc_vec[1]~q ;
wire \wd_vec[1]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][1]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][1]~q ;
wire \delay_ctrl_np|tdl_arr[9]~q ;
wire \wc_vec[0]~q ;
wire \wd_vec[0]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][0][0]~q ;
wire \gen_dft_1:bfpdft|reg_no_twiddle[6][1][0]~q ;
wire \twiddle_data[0][1][0]~q ;
wire \twiddle_data[0][1][1]~q ;
wire \twiddle_data[0][1][2]~q ;
wire \twiddle_data[0][1][3]~q ;
wire \twiddle_data[0][1][4]~q ;
wire \twiddle_data[0][1][5]~q ;
wire \twiddle_data[0][1][6]~q ;
wire \twiddle_data[0][1][7]~q ;
wire \twiddle_data[0][0][7]~q ;
wire \twiddle_data[1][0][7]~q ;
wire \twiddle_data[1][1][0]~q ;
wire \twiddle_data[1][1][1]~q ;
wire \twiddle_data[1][1][2]~q ;
wire \twiddle_data[1][1][3]~q ;
wire \twiddle_data[1][1][4]~q ;
wire \twiddle_data[1][1][5]~q ;
wire \twiddle_data[1][1][6]~q ;
wire \twiddle_data[1][1][7]~q ;
wire \twiddle_data[2][0][7]~q ;
wire \twiddle_data[2][1][0]~q ;
wire \twiddle_data[2][1][1]~q ;
wire \twiddle_data[2][1][2]~q ;
wire \twiddle_data[2][1][3]~q ;
wire \twiddle_data[2][1][4]~q ;
wire \twiddle_data[2][1][5]~q ;
wire \twiddle_data[2][1][6]~q ;
wire \twiddle_data[2][1][7]~q ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \data_rdy_vec[10]~q ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \data_rdy_vec[9]~q ;
wire \wren_b[1]~q ;
wire \ccc|b_ram_data_in_bus[46]~q ;
wire \ccc|wraddress_b_bus[0]~q ;
wire \ccc|wraddress_b_bus[9]~q ;
wire \ccc|wraddress_b_bus[10]~q ;
wire \ccc|wraddress_b_bus[11]~q ;
wire \ccc|rdaddress_b_bus[0]~q ;
wire \ccc|rdaddress_b_bus[9]~q ;
wire \ccc|rdaddress_b_bus[10]~q ;
wire \ccc|rdaddress_b_bus[11]~q ;
wire \wren_a[1]~q ;
wire \ccc|a_ram_data_in_bus[46]~q ;
wire \ccc|wraddress_a_bus[0]~q ;
wire \ccc|wraddress_a_bus[9]~q ;
wire \ccc|wraddress_a_bus[10]~q ;
wire \ccc|wraddress_a_bus[11]~q ;
wire \ccc|rdaddress_a_bus[0]~q ;
wire \ccc|rdaddress_a_bus[9]~q ;
wire \ccc|rdaddress_a_bus[10]~q ;
wire \ccc|rdaddress_a_bus[11]~q ;
wire \wren_b[2]~q ;
wire \ccc|b_ram_data_in_bus[30]~q ;
wire \ccc|wraddress_b_bus[12]~q ;
wire \ccc|wraddress_b_bus[5]~q ;
wire \ccc|rdaddress_b_bus[12]~q ;
wire \ccc|rdaddress_b_bus[5]~q ;
wire \wren_a[2]~q ;
wire \ccc|a_ram_data_in_bus[30]~q ;
wire \ccc|wraddress_a_bus[12]~q ;
wire \ccc|wraddress_a_bus[5]~q ;
wire \ccc|rdaddress_a_bus[12]~q ;
wire \ccc|rdaddress_a_bus[5]~q ;
wire \wren_b[3]~q ;
wire \ccc|b_ram_data_in_bus[14]~q ;
wire \ccc|wraddress_b_bus[1]~q ;
wire \ccc|rdaddress_b_bus[1]~q ;
wire \wren_a[3]~q ;
wire \ccc|a_ram_data_in_bus[14]~q ;
wire \ccc|wraddress_a_bus[1]~q ;
wire \ccc|rdaddress_a_bus[1]~q ;
wire \wren_b[0]~q ;
wire \ccc|b_ram_data_in_bus[62]~q ;
wire \ccc|wraddress_b_bus[13]~q ;
wire \ccc|rdaddress_b_bus[13]~q ;
wire \wren_a[0]~q ;
wire \ccc|a_ram_data_in_bus[62]~q ;
wire \ccc|wraddress_a_bus[13]~q ;
wire \ccc|rdaddress_a_bus[13]~q ;
wire \ccc|b_ram_data_in_bus[45]~q ;
wire \ccc|a_ram_data_in_bus[45]~q ;
wire \ccc|b_ram_data_in_bus[29]~q ;
wire \ccc|a_ram_data_in_bus[29]~q ;
wire \ccc|b_ram_data_in_bus[13]~q ;
wire \ccc|a_ram_data_in_bus[13]~q ;
wire \ccc|b_ram_data_in_bus[61]~q ;
wire \ccc|a_ram_data_in_bus[61]~q ;
wire \ccc|b_ram_data_in_bus[42]~q ;
wire \ccc|a_ram_data_in_bus[42]~q ;
wire \ccc|b_ram_data_in_bus[26]~q ;
wire \ccc|a_ram_data_in_bus[26]~q ;
wire \ccc|b_ram_data_in_bus[10]~q ;
wire \ccc|a_ram_data_in_bus[10]~q ;
wire \ccc|b_ram_data_in_bus[58]~q ;
wire \ccc|a_ram_data_in_bus[58]~q ;
wire \ccc|b_ram_data_in_bus[43]~q ;
wire \ccc|a_ram_data_in_bus[43]~q ;
wire \ccc|b_ram_data_in_bus[27]~q ;
wire \ccc|a_ram_data_in_bus[27]~q ;
wire \ccc|b_ram_data_in_bus[11]~q ;
wire \ccc|a_ram_data_in_bus[11]~q ;
wire \ccc|b_ram_data_in_bus[59]~q ;
wire \ccc|a_ram_data_in_bus[59]~q ;
wire \ccc|b_ram_data_in_bus[44]~q ;
wire \ccc|a_ram_data_in_bus[44]~q ;
wire \ccc|b_ram_data_in_bus[28]~q ;
wire \ccc|a_ram_data_in_bus[28]~q ;
wire \ccc|b_ram_data_in_bus[12]~q ;
wire \ccc|a_ram_data_in_bus[12]~q ;
wire \ccc|b_ram_data_in_bus[60]~q ;
wire \ccc|a_ram_data_in_bus[60]~q ;
wire \ccc|b_ram_data_in_bus[47]~q ;
wire \ccc|a_ram_data_in_bus[47]~q ;
wire \ccc|b_ram_data_in_bus[31]~q ;
wire \ccc|a_ram_data_in_bus[31]~q ;
wire \ccc|b_ram_data_in_bus[15]~q ;
wire \ccc|a_ram_data_in_bus[15]~q ;
wire \ccc|b_ram_data_in_bus[63]~q ;
wire \ccc|a_ram_data_in_bus[63]~q ;
wire \ccc|b_ram_data_in_bus[39]~q ;
wire \ccc|a_ram_data_in_bus[39]~q ;
wire \ccc|b_ram_data_in_bus[23]~q ;
wire \ccc|a_ram_data_in_bus[23]~q ;
wire \ccc|b_ram_data_in_bus[7]~q ;
wire \ccc|a_ram_data_in_bus[7]~q ;
wire \ccc|b_ram_data_in_bus[55]~q ;
wire \ccc|a_ram_data_in_bus[55]~q ;
wire \ccc|b_ram_data_in_bus[38]~q ;
wire \ccc|a_ram_data_in_bus[38]~q ;
wire \ccc|b_ram_data_in_bus[22]~q ;
wire \ccc|a_ram_data_in_bus[22]~q ;
wire \ccc|b_ram_data_in_bus[6]~q ;
wire \ccc|a_ram_data_in_bus[6]~q ;
wire \ccc|b_ram_data_in_bus[54]~q ;
wire \ccc|a_ram_data_in_bus[54]~q ;
wire \ccc|b_ram_data_in_bus[35]~q ;
wire \ccc|a_ram_data_in_bus[35]~q ;
wire \ccc|b_ram_data_in_bus[19]~q ;
wire \ccc|a_ram_data_in_bus[19]~q ;
wire \ccc|b_ram_data_in_bus[3]~q ;
wire \ccc|a_ram_data_in_bus[3]~q ;
wire \ccc|b_ram_data_in_bus[51]~q ;
wire \ccc|a_ram_data_in_bus[51]~q ;
wire \ccc|b_ram_data_in_bus[36]~q ;
wire \ccc|a_ram_data_in_bus[36]~q ;
wire \ccc|b_ram_data_in_bus[20]~q ;
wire \ccc|a_ram_data_in_bus[20]~q ;
wire \ccc|b_ram_data_in_bus[4]~q ;
wire \ccc|a_ram_data_in_bus[4]~q ;
wire \ccc|b_ram_data_in_bus[52]~q ;
wire \ccc|a_ram_data_in_bus[52]~q ;
wire \ccc|b_ram_data_in_bus[37]~q ;
wire \ccc|a_ram_data_in_bus[37]~q ;
wire \ccc|b_ram_data_in_bus[21]~q ;
wire \ccc|a_ram_data_in_bus[21]~q ;
wire \ccc|b_ram_data_in_bus[5]~q ;
wire \ccc|a_ram_data_in_bus[5]~q ;
wire \ccc|b_ram_data_in_bus[53]~q ;
wire \ccc|a_ram_data_in_bus[53]~q ;
wire \ccc|b_ram_data_in_bus[34]~q ;
wire \ccc|a_ram_data_in_bus[34]~q ;
wire \ccc|b_ram_data_in_bus[18]~q ;
wire \ccc|a_ram_data_in_bus[18]~q ;
wire \ccc|b_ram_data_in_bus[2]~q ;
wire \ccc|a_ram_data_in_bus[2]~q ;
wire \ccc|b_ram_data_in_bus[50]~q ;
wire \ccc|a_ram_data_in_bus[50]~q ;
wire \ccc|b_ram_data_in_bus[24]~q ;
wire \ccc|a_ram_data_in_bus[24]~q ;
wire \ccc|b_ram_data_in_bus[8]~q ;
wire \ccc|a_ram_data_in_bus[8]~q ;
wire \ccc|b_ram_data_in_bus[56]~q ;
wire \ccc|a_ram_data_in_bus[56]~q ;
wire \ccc|b_ram_data_in_bus[40]~q ;
wire \ccc|a_ram_data_in_bus[40]~q ;
wire \ccc|b_ram_data_in_bus[25]~q ;
wire \ccc|a_ram_data_in_bus[25]~q ;
wire \ccc|b_ram_data_in_bus[9]~q ;
wire \ccc|a_ram_data_in_bus[9]~q ;
wire \ccc|b_ram_data_in_bus[57]~q ;
wire \ccc|a_ram_data_in_bus[57]~q ;
wire \ccc|b_ram_data_in_bus[41]~q ;
wire \ccc|a_ram_data_in_bus[41]~q ;
wire \ccc|b_ram_data_in_bus[0]~q ;
wire \ccc|a_ram_data_in_bus[0]~q ;
wire \ccc|b_ram_data_in_bus[48]~q ;
wire \ccc|a_ram_data_in_bus[48]~q ;
wire \ccc|b_ram_data_in_bus[32]~q ;
wire \ccc|a_ram_data_in_bus[32]~q ;
wire \ccc|b_ram_data_in_bus[16]~q ;
wire \ccc|a_ram_data_in_bus[16]~q ;
wire \ccc|b_ram_data_in_bus[1]~q ;
wire \ccc|a_ram_data_in_bus[1]~q ;
wire \ccc|b_ram_data_in_bus[49]~q ;
wire \ccc|a_ram_data_in_bus[49]~q ;
wire \ccc|b_ram_data_in_bus[33]~q ;
wire \ccc|a_ram_data_in_bus[33]~q ;
wire \ccc|b_ram_data_in_bus[17]~q ;
wire \ccc|a_ram_data_in_bus[17]~q ;
wire \data_rdy_vec[8]~q ;
wire \writer|wren[1]~q ;
wire \writer|data_in_r[6]~q ;
wire \writer|wr_address_i_int[0]~q ;
wire \writer|wr_address_i_int[1]~q ;
wire \writer|wr_address_i_int[2]~q ;
wire \writer|wr_address_i_int[3]~q ;
wire \writer|wren[2]~q ;
wire \writer|wren[3]~q ;
wire \writer|wren[0]~q ;
wire \writer|data_in_r[5]~q ;
wire \writer|data_in_r[2]~q ;
wire \writer|data_in_r[3]~q ;
wire \writer|data_in_r[4]~q ;
wire \writer|data_in_r[7]~q ;
wire \writer|data_in_i[7]~q ;
wire \writer|data_in_i[6]~q ;
wire \writer|data_in_i[3]~q ;
wire \writer|data_in_i[4]~q ;
wire \writer|data_in_i[5]~q ;
wire \writer|data_in_i[2]~q ;
wire \writer|data_in_r[0]~q ;
wire \writer|data_in_r[1]~q ;
wire \writer|data_in_i[0]~q ;
wire \writer|data_in_i[1]~q ;
wire \data_rdy_vec[7]~q ;
wire \core_real_in[6]~q ;
wire \core_real_in[5]~q ;
wire \core_real_in[2]~q ;
wire \core_real_in[3]~q ;
wire \core_real_in[4]~q ;
wire \core_real_in[7]~q ;
wire \core_imag_in[7]~q ;
wire \core_imag_in[6]~q ;
wire \core_imag_in[3]~q ;
wire \core_imag_in[4]~q ;
wire \core_imag_in[5]~q ;
wire \core_imag_in[2]~q ;
wire \core_real_in[0]~q ;
wire \core_real_in[1]~q ;
wire \core_imag_in[0]~q ;
wire \core_imag_in[1]~q ;
wire \data_rdy_vec[6]~q ;
wire \writer|anb~q ;
wire \data_real_in_reg[6]~q ;
wire \data_imag_in_reg[6]~q ;
wire \data_real_in_reg[5]~q ;
wire \data_imag_in_reg[5]~q ;
wire \data_real_in_reg[2]~q ;
wire \data_imag_in_reg[2]~q ;
wire \data_real_in_reg[3]~q ;
wire \data_imag_in_reg[3]~q ;
wire \data_real_in_reg[4]~q ;
wire \data_imag_in_reg[4]~q ;
wire \data_real_in_reg[7]~q ;
wire \data_imag_in_reg[7]~q ;
wire \data_real_in_reg[0]~q ;
wire \data_imag_in_reg[0]~q ;
wire \data_real_in_reg[1]~q ;
wire \data_imag_in_reg[1]~q ;
wire \data_rdy_vec[5]~q ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \data_count_sig[2]~5_combout ;
wire \auk_dsp_interface_controller_1|source_packet_error[1]~q ;
wire \auk_dsp_interface_controller_1|source_packet_error[0]~q ;
wire \auk_dsp_atlantic_sink_1|sink_stall~combout ;
wire \auk_dsp_interface_controller_1|sink_stall_reg~q ;
wire \auk_dsp_interface_controller_1|source_stall_reg~q ;
wire \auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ;
wire \master_sink_ena~q ;
wire \auk_dsp_atlantic_sink_1|send_eop_s~q ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[1]~q ;
wire \auk_dsp_atlantic_sink_1|packet_error_s[0]~q ;
wire \sink_ready_ctrl_d~q ;
wire \auk_dsp_atlantic_sink_1|send_sop_s~q ;
wire \sop~q ;
wire \auk_dsp_atlantic_source_1|stall_controller_comb~0_combout ;
wire \data_count_sig[3]~q ;
wire \data_count_sig[2]~q ;
wire \data_count_sig[1]~q ;
wire \data_count_sig[0]~q ;
wire \data_count_sig[5]~q ;
wire \auk_dsp_atlantic_source_1|source_stall_int_d~q ;
wire \auk_dsp_interface_controller_1|stall_reg~q ;
wire \data_count_sig[4]~q ;
wire \exponent_out[0]~q ;
wire \exponent_out[1]~q ;
wire \exponent_out[2]~q ;
wire \exponent_out[3]~q ;
wire \exponent_out[4]~q ;
wire \exponent_out[5]~q ;
wire \auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ;
wire \auk_dsp_atlantic_source_1|Mux0~0_combout ;
wire \auk_dsp_atlantic_source_1|Mux0~1_combout ;
wire \auk_dsp_atlantic_source_1|Mux0~2_combout ;
wire \global_clock_enable~0_combout ;
wire \sink_in_work~0_combout ;
wire \sop~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \data_sample_counter~0_combout ;
wire \master_source_sop~q ;
wire \data_count_sig[3]~0_combout ;
wire \data_count_sig[1]~1_combout ;
wire \data_count_sig~2_combout ;
wire \LessThan0~2_combout ;
wire \data_count_sig[5]~3_combout ;
wire \auk_dsp_atlantic_source_1|stall_controller_comb~1_combout ;
wire \data_count_sig[4]~4_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[0]~q ;
wire \fft_imag_out[1]~0_combout ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[1]~q ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[2]~q ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[3]~q ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[4]~q ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[5]~q ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[6]~q ;
wire \gen_radix_4_last_pass:lpp|data_imag_o[7]~q ;
wire \blk_exp_accum[0]~q ;
wire \exponent_out~0_combout ;
wire \blk_exp_accum[1]~q ;
wire \exponent_out~1_combout ;
wire \blk_exp_accum[2]~q ;
wire \exponent_out~2_combout ;
wire \blk_exp_accum[3]~q ;
wire \exponent_out~3_combout ;
wire \blk_exp_accum[4]~q ;
wire \exponent_out~4_combout ;
wire \blk_exp_accum[5]~q ;
wire \exponent_out~5_combout ;
wire \fft_s2_cur.IDLE~q ;
wire \WideNor1~combout ;
wire \master_source_sop~0_combout ;
wire \fft_s2_cur.FIRST_LPP_C~q ;
wire \fft_dirn_stream~0_combout ;
wire \gen_dft_1:bfpc|blk_exp[0]~q ;
wire \Selector5~0_combout ;
wire \gen_dft_1:bfpc|blk_exp[1]~q ;
wire \Selector4~0_combout ;
wire \gen_dft_1:bfpc|blk_exp[2]~q ;
wire \Selector3~0_combout ;
wire \gen_dft_1:bfpc|blk_exp[3]~q ;
wire \Selector2~0_combout ;
wire \gen_dft_1:bfpc|blk_exp[4]~q ;
wire \Selector1~0_combout ;
wire \gen_dft_1:bfpc|blk_exp[5]~q ;
wire \Selector0~0_combout ;
wire \fft_s2_cur.LPP_C_OUTPUT~q ;
wire \lpp_count_offset[0]~q ;
wire \fft_s2_cur.IDLE~0_combout ;
wire \fft_s2_cur.IDLE~1_combout ;
wire \fft_s2_cur.LAST_LPP_C~q ;
wire \Selector17~0_combout ;
wire \fft_dirn_held_o2~0_combout ;
wire \fft_s2_cur~9_combout ;
wire \fft_s2_cur.LPP_C_OUTPUT~0_combout ;
wire \Add1~0_combout ;
wire \lpp_count_offset[0]~0_combout ;
wire \lpp_count_offset~1_combout ;
wire \Add1~1_combout ;
wire \Add1~2_combout ;
wire \Add1~3_combout ;
wire \Add1~4_combout ;
wire \fft_s2_cur.LAST_LPP_C~0_combout ;
wire \fft_dirn_held_o~0_combout ;
wire \gen_le256_mk:ctrl|p[1]~q ;
wire \Selector11~0_combout ;
wire \Selector10~0_combout ;
wire \lpp_count~0_combout ;
wire \Selector9~0_combout ;
wire \Selector8~0_combout ;
wire \Selector7~0_combout ;
wire \gen_dft_1:bfpc|slb_last[0]~q ;
wire \gen_dft_1:bfpc|slb_last[1]~q ;
wire \gen_dft_1:bfpc|slb_last[2]~q ;
wire \inv_i~q ;
wire \fft_dirn~0_combout ;
wire \gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[0]~q ;
wire \gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[1]~q ;
wire \gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[2]~q ;
wire \inv_i~0_combout ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][4]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][4]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][4]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][4]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][4]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][4]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][5]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][5]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][5]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][5]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][5]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][5]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][6]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][6]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][6]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][6]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][6]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][2]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][3]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][4]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][5]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][6]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][7]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][1]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][1]~q ;
wire \lpp_ram_data_out~0_combout ;
wire \lpp_ram_data_out~1_combout ;
wire \lpp_ram_data_out~2_combout ;
wire \lpp_ram_data_out~3_combout ;
wire \lpp_ram_data_out~4_combout ;
wire \lpp_ram_data_out~5_combout ;
wire \lpp_ram_data_out~6_combout ;
wire \lpp_ram_data_out~7_combout ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][0]~q ;
wire \gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][0]~q ;
wire \lpp_ram_data_out~8_combout ;
wire \lpp_ram_data_out~9_combout ;
wire \lpp_ram_data_out~10_combout ;
wire \lpp_ram_data_out~11_combout ;
wire \lpp_ram_data_out~12_combout ;
wire \lpp_ram_data_out~13_combout ;
wire \lpp_ram_data_out~14_combout ;
wire \lpp_ram_data_out~15_combout ;
wire \lpp_ram_data_out~16_combout ;
wire \lpp_ram_data_out~17_combout ;
wire \lpp_ram_data_out~18_combout ;
wire \lpp_ram_data_out~19_combout ;
wire \lpp_ram_data_out~20_combout ;
wire \lpp_ram_data_out~21_combout ;
wire \lpp_ram_data_out~22_combout ;
wire \lpp_ram_data_out~23_combout ;
wire \lpp_ram_data_out~24_combout ;
wire \lpp_ram_data_out~25_combout ;
wire \lpp_ram_data_out~26_combout ;
wire \lpp_ram_data_out~27_combout ;
wire \lpp_ram_data_out~28_combout ;
wire \lpp_ram_data_out~29_combout ;
wire \lpp_ram_data_out~30_combout ;
wire \lpp_ram_data_out~31_combout ;
wire \lpp_ram_data_out~32_combout ;
wire \lpp_ram_data_out~33_combout ;
wire \lpp_ram_data_out~34_combout ;
wire \lpp_ram_data_out~35_combout ;
wire \lpp_ram_data_out~36_combout ;
wire \lpp_ram_data_out~37_combout ;
wire \lpp_ram_data_out~38_combout ;
wire \lpp_ram_data_out~39_combout ;
wire \lpp_ram_data_out~40_combout ;
wire \lpp_ram_data_out~41_combout ;
wire \lpp_ram_data_out~42_combout ;
wire \lpp_ram_data_out~43_combout ;
wire \lpp_ram_data_out~44_combout ;
wire \lpp_ram_data_out~45_combout ;
wire \lpp_ram_data_out~46_combout ;
wire \lpp_ram_data_out~47_combout ;
wire \ram_cxb_wr_data|ram_in_reg[3][2]~q ;
wire \gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][0]~q ;
wire \gen_wrsw_1:ram_cxb_wr|ram_in_reg[3][1]~q ;
wire \lpp_sel~0_combout ;
wire \ram_cxb_wr_data|ram_in_reg[0][2]~q ;
wire \gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][0]~q ;
wire \gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][2]~q ;
wire \gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][2]~q ;
wire \gen_wrsw_1:ram_cxb_wr|ram_in_reg[2][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][2]~q ;
wire \lpp_ram_data_out~48_combout ;
wire \lpp_ram_data_out~49_combout ;
wire \lpp_ram_data_out~50_combout ;
wire \lpp_ram_data_out~51_combout ;
wire \lpp_ram_data_out~52_combout ;
wire \lpp_ram_data_out~53_combout ;
wire \lpp_ram_data_out~54_combout ;
wire \lpp_ram_data_out~55_combout ;
wire \ram_cxb_wr_data|ram_in_reg[3][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][3]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][4]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][5]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][6]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][7]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][7]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][2]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][2]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][2]~q ;
wire \ram_cxb_rd|ram_in_reg[0][2]~q ;
wire \ram_cxb_rd|ram_in_reg[0][3]~q ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[1][2]~q ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[3][3]~q ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][2]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][2]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][2]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][1]~q ;
wire \lpp_ram_data_out~56_combout ;
wire \lpp_ram_data_out~57_combout ;
wire \lpp_ram_data_out~58_combout ;
wire \lpp_ram_data_out~59_combout ;
wire \lpp_ram_data_out~60_combout ;
wire \lpp_ram_data_out~61_combout ;
wire \lpp_ram_data_out~62_combout ;
wire \lpp_ram_data_out~63_combout ;
wire \en_slb~q ;
wire \p_tdl[0][0]~q ;
wire \p_tdl[0][1]~q ;
wire \gen_le256_mk:ctrl|k_count[1]~q ;
wire \gen_le256_mk:ctrl|k_count[3]~q ;
wire \gen_le256_mk:ctrl|k_count[0]~q ;
wire \gen_le256_mk:ctrl|k_count[2]~q ;
wire \ram_cxb_rd|ram_in_reg[0][0]~q ;
wire \ram_cxb_rd|ram_in_reg[1][0]~q ;
wire \ram_cxb_rd|ram_in_reg[3][1]~q ;
wire \ram_cxb_rd|ram_in_reg[1][1]~q ;
wire \ram_cxb_rd|ram_in_reg[2][1]~q ;
wire \ram_cxb_rd|ram_in_reg[0][1]~q ;
wire \rd_adgen|rd_addr_d[2]~q ;
wire \rd_adgen|rd_addr_d[3]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[0]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[1]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|sw[0]~q ;
wire \gen_radix_4_last_pass:gen_lpp_addr|sw[1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][1]~q ;
wire \ram_cxb_wr_data|ram_in_reg[3][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[0][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[1][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[2][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[7][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[4][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[5][0]~q ;
wire \ram_cxb_wr_data|ram_in_reg[6][0]~q ;
wire \en_slb~0_combout ;
wire \rd_adgen|rd_addr_d[0]~q ;
wire \rd_adgen|sw[0]~q ;
wire \rd_adgen|rd_addr_c[0]~q ;
wire \rd_adgen|rd_addr_b[1]~q ;
wire \rd_adgen|sw[1]~q ;
wire \rd_adgen|rd_addr_d[1]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][0]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][0]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][0]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][0]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][0]~q ;
wire \gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][0]~q ;
wire \sel_we|wc_i~q ;
wire \sel_we|wd_i~q ;
wire \ram_a_not_b_vec[26]~q ;
wire \p_cd_en[0]~q ;
wire \p_cd_en[1]~q ;
wire \twiddle_data[0][0][0]~q ;
wire \twiddle_data[0][0][1]~q ;
wire \twiddle_data[0][0][2]~q ;
wire \twiddle_data[0][0][3]~q ;
wire \twiddle_data[0][0][4]~q ;
wire \twiddle_data[0][0][5]~q ;
wire \twiddle_data[0][0][6]~q ;
wire \twiddle_data[1][0][0]~q ;
wire \twiddle_data[1][0][1]~q ;
wire \twiddle_data[1][0][2]~q ;
wire \twiddle_data[1][0][3]~q ;
wire \twiddle_data[1][0][4]~q ;
wire \twiddle_data[1][0][5]~q ;
wire \twiddle_data[1][0][6]~q ;
wire \twiddle_data[2][0][0]~q ;
wire \twiddle_data[2][0][1]~q ;
wire \twiddle_data[2][0][2]~q ;
wire \twiddle_data[2][0][3]~q ;
wire \twiddle_data[2][0][4]~q ;
wire \twiddle_data[2][0][5]~q ;
wire \twiddle_data[2][0][6]~q ;
wire \ram_a_not_b_vec[25]~q ;
wire \ram_a_not_b_vec~0_combout ;
wire \p_tdl[12][0]~q ;
wire \p_tdl[12][1]~q ;
wire \twiddle_data~0_combout ;
wire \twiddle_data~1_combout ;
wire \twiddle_data~2_combout ;
wire \twiddle_data~3_combout ;
wire \twiddle_data~4_combout ;
wire \twiddle_data~5_combout ;
wire \twiddle_data~6_combout ;
wire \twiddle_data~7_combout ;
wire \twiddle_data~8_combout ;
wire \twiddle_data~9_combout ;
wire \twiddle_data~10_combout ;
wire \twiddle_data~11_combout ;
wire \twiddle_data~12_combout ;
wire \twiddle_data~13_combout ;
wire \twiddle_data~14_combout ;
wire \twiddle_data~15_combout ;
wire \twiddle_data~16_combout ;
wire \twiddle_data~17_combout ;
wire \twiddle_data~18_combout ;
wire \twiddle_data~19_combout ;
wire \twiddle_data~20_combout ;
wire \ram_a_not_b_vec[24]~q ;
wire \ram_a_not_b_vec~1_combout ;
wire \p_tdl[11][0]~q ;
wire \p_tdl[11][1]~q ;
wire \twid_factors|twad_tdl[6][0]~q ;
wire \twid_factors|twad_tdl[6][1]~q ;
wire \twid_factors|twad_tdl[6][2]~q ;
wire \twid_factors|twad_tdl[6][3]~q ;
wire \ram_a_not_b_vec[23]~q ;
wire \ram_a_not_b_vec~2_combout ;
wire \p_tdl[10][0]~q ;
wire \p_tdl[10][1]~q ;
wire \ram_a_not_b_vec[22]~q ;
wire \ram_a_not_b_vec~3_combout ;
wire \p_tdl[9][0]~q ;
wire \p_tdl[9][1]~q ;
wire \ram_a_not_b_vec[21]~q ;
wire \ram_a_not_b_vec~4_combout ;
wire \p_tdl[8][0]~q ;
wire \p_tdl[8][1]~q ;
wire \ram_a_not_b_vec[20]~q ;
wire \ram_a_not_b_vec~5_combout ;
wire \p_tdl[7][0]~q ;
wire \p_tdl[7][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][7]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][6]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][3]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][4]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][5]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][2]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][2]~q ;
wire \ram_a_not_b_vec[19]~q ;
wire \ram_a_not_b_vec~6_combout ;
wire \p_tdl[6][0]~q ;
wire \p_tdl[6][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[2][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[0][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[7][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[5][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[3][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[1][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[6][1]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][0]~q ;
wire \ram_cxb_bfp_data|ram_in_reg[4][1]~q ;
wire \ccc|ram_data_out1[14]~q ;
wire \ccc|ram_data_out2[14]~q ;
wire \ccc|ram_data_out3[14]~q ;
wire \ccc|ram_data_out0[14]~q ;
wire \sw_r_tdl[4][0]~q ;
wire \sw_r_tdl[4][1]~q ;
wire \ccc|ram_data_out1[13]~q ;
wire \ccc|ram_data_out2[13]~q ;
wire \ccc|ram_data_out3[13]~q ;
wire \ccc|ram_data_out0[13]~q ;
wire \ccc|ram_data_out1[10]~q ;
wire \ccc|ram_data_out2[10]~q ;
wire \ccc|ram_data_out3[10]~q ;
wire \ccc|ram_data_out0[10]~q ;
wire \ccc|ram_data_out1[11]~q ;
wire \ccc|ram_data_out2[11]~q ;
wire \ccc|ram_data_out3[11]~q ;
wire \ccc|ram_data_out0[11]~q ;
wire \ccc|ram_data_out1[12]~q ;
wire \ccc|ram_data_out2[12]~q ;
wire \ccc|ram_data_out3[12]~q ;
wire \ccc|ram_data_out0[12]~q ;
wire \ccc|ram_data_out1[15]~q ;
wire \ccc|ram_data_out2[15]~q ;
wire \ccc|ram_data_out3[15]~q ;
wire \ccc|ram_data_out0[15]~q ;
wire \ccc|ram_data_out1[7]~q ;
wire \ccc|ram_data_out2[7]~q ;
wire \ccc|ram_data_out3[7]~q ;
wire \ccc|ram_data_out0[7]~q ;
wire \ccc|ram_data_out1[6]~q ;
wire \ccc|ram_data_out2[6]~q ;
wire \ccc|ram_data_out3[6]~q ;
wire \ccc|ram_data_out0[6]~q ;
wire \ccc|ram_data_out1[3]~q ;
wire \ccc|ram_data_out2[3]~q ;
wire \ccc|ram_data_out3[3]~q ;
wire \ccc|ram_data_out0[3]~q ;
wire \ccc|ram_data_out1[4]~q ;
wire \ccc|ram_data_out2[4]~q ;
wire \ccc|ram_data_out3[4]~q ;
wire \ccc|ram_data_out0[4]~q ;
wire \ccc|ram_data_out1[5]~q ;
wire \ccc|ram_data_out2[5]~q ;
wire \ccc|ram_data_out3[5]~q ;
wire \ccc|ram_data_out0[5]~q ;
wire \ccc|ram_data_out1[2]~q ;
wire \ccc|ram_data_out2[2]~q ;
wire \ccc|ram_data_out3[2]~q ;
wire \ccc|ram_data_out0[2]~q ;
wire \ram_a_not_b_vec[18]~q ;
wire \ram_a_not_b_vec~7_combout ;
wire \p_tdl[5][0]~q ;
wire \p_tdl[5][1]~q ;
wire \ccc|ram_data_out2[8]~q ;
wire \ccc|ram_data_out3[8]~q ;
wire \ccc|ram_data_out0[8]~q ;
wire \ccc|ram_data_out1[8]~q ;
wire \ccc|ram_data_out2[9]~q ;
wire \ccc|ram_data_out3[9]~q ;
wire \ccc|ram_data_out0[9]~q ;
wire \ccc|ram_data_out1[9]~q ;
wire \ccc|ram_data_out3[0]~q ;
wire \ccc|ram_data_out0[0]~q ;
wire \ccc|ram_data_out1[0]~q ;
wire \ccc|ram_data_out2[0]~q ;
wire \ccc|ram_data_out3[1]~q ;
wire \ccc|ram_data_out0[1]~q ;
wire \ccc|ram_data_out1[1]~q ;
wire \ccc|ram_data_out2[1]~q ;
wire \ram_a_not_b_vec[10]~q ;
wire \sw_r_tdl[3][0]~q ;
wire \sw_r_tdl[3][1]~q ;
wire \ram_a_not_b_vec[17]~q ;
wire \ram_a_not_b_vec~8_combout ;
wire \p_tdl[4][0]~q ;
wire \p_tdl[4][1]~q ;
wire \ram_a_not_b_vec[9]~q ;
wire \ram_a_not_b_vec~9_combout ;
wire \sw_r_tdl[2][0]~q ;
wire \sw_r_tdl[2][1]~q ;
wire \ram_a_not_b_vec[16]~q ;
wire \ram_a_not_b_vec~10_combout ;
wire \p_tdl[3][0]~q ;
wire \p_tdl[3][1]~q ;
wire \rd_adgen|Mux1~1_combout ;
wire \rd_adgen|Mux0~1_combout ;
wire \rd_adgen|Mux1~2_combout ;
wire \rd_adgen|Mux0~2_combout ;
wire \ram_a_not_b_vec[8]~q ;
wire \ram_a_not_b_vec~11_combout ;
wire \ram_a_not_b_vec[1]~q ;
wire \wren_b~0_combout ;
wire \ram_a_not_b_vec[7]~q ;
wire \sel_anb_addr~combout ;
wire \wren_a~0_combout ;
wire \wren_b~1_combout ;
wire \wren_a~1_combout ;
wire \wren_b~2_combout ;
wire \wren_a~2_combout ;
wire \wren_b~3_combout ;
wire \wren_a~3_combout ;
wire \sw_r_tdl[1][0]~q ;
wire \sw_r_tdl[1][1]~q ;
wire \ram_a_not_b_vec[15]~q ;
wire \ram_a_not_b_vec~12_combout ;
wire \p_tdl[2][0]~q ;
wire \p_tdl[2][1]~q ;
wire \ram_a_not_b_vec~13_combout ;
wire \ram_a_not_b_vec[0]~q ;
wire \ram_a_not_b_vec~14_combout ;
wire \ram_a_not_b_vec[6]~q ;
wire \ram_a_not_b_vec~15_combout ;
wire \sw_r_tdl[0][0]~q ;
wire \sw_r_tdl[0][1]~q ;
wire \ram_a_not_b_vec[14]~q ;
wire \ram_a_not_b_vec~16_combout ;
wire \p_tdl[1][0]~q ;
wire \p_tdl[1][1]~q ;
wire \ram_a_not_b_vec~17_combout ;
wire \ram_a_not_b_vec[5]~q ;
wire \ram_a_not_b_vec~18_combout ;
wire \ram_a_not_b_vec[13]~q ;
wire \ram_a_not_b_vec~19_combout ;
wire \ram_a_not_b_vec[4]~q ;
wire \ram_a_not_b_vec~20_combout ;
wire \ram_a_not_b_vec[12]~q ;
wire \ram_a_not_b_vec~21_combout ;
wire \ram_a_not_b_vec[3]~q ;
wire \ram_a_not_b_vec~22_combout ;
wire \ram_a_not_b_vec[11]~q ;
wire \ram_a_not_b_vec~23_combout ;
wire \ram_a_not_b_vec[2]~q ;
wire \ram_a_not_b_vec~24_combout ;
wire \ram_a_not_b_vec~25_combout ;
wire \ram_a_not_b_vec~26_combout ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][3]~_wirecell_combout ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[1][2]~_wirecell_combout ;
wire \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[3][3]~_wirecell_combout ;


IFFT_auk_dspip_avalon_streaming_sink auk_dsp_atlantic_sink_1(
	.sink_in_work(\sink_in_work~q ),
	.q_b_14(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_6(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_13(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_5(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_10(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_2(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_11(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_3(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_12(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_4(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_15(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_7(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_8(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_0(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_9(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_1(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.at_sink_ready_s1(at_sink_ready_s),
	.sink_stall1(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.sink_stall_reg(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.source_stall_reg(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.master_sink_ena(\master_sink_ena~q ),
	.send_eop_s1(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.send_sop_s1(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.sink_ready_ctrl1(\auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.sink_eop(sink_eop),
	.sink_valid(sink_valid),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.sink_sop(sink_sop),
	.at_sink_data({sink_real[7],sink_real[6],sink_real[5],sink_real[4],sink_real[3],sink_real[2],sink_real[1],sink_real[0],sink_imag[7],sink_imag[6],sink_imag[5],sink_imag[4],sink_imag[3],sink_imag[2],sink_imag[1],sink_imag[0]}));

IFFT_asj_fft_dft_bfp \gen_dft_1:bfpdft (
	.next_block(\writer|next_block~q ),
	.reg_no_twiddle603(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][3]~q ),
	.reg_no_twiddle607(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][7]~q ),
	.reg_no_twiddle617(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][7]~q ),
	.reg_no_twiddle613(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][3]~q ),
	.reg_no_twiddle604(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][4]~q ),
	.reg_no_twiddle614(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][4]~q ),
	.reg_no_twiddle605(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][5]~q ),
	.reg_no_twiddle615(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][5]~q ),
	.reg_no_twiddle606(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][6]~q ),
	.reg_no_twiddle616(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][6]~q ),
	.reg_no_twiddle602(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][2]~q ),
	.reg_no_twiddle612(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][2]~q ),
	.reg_no_twiddle601(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][1]~q ),
	.reg_no_twiddle611(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][1]~q ),
	.tdl_arr_9(\delay_ctrl_np|tdl_arr[9]~q ),
	.reg_no_twiddle600(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][0]~q ),
	.reg_no_twiddle610(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][0]~q ),
	.twiddle_data010(\twiddle_data[0][1][0]~q ),
	.twiddle_data011(\twiddle_data[0][1][1]~q ),
	.twiddle_data012(\twiddle_data[0][1][2]~q ),
	.twiddle_data013(\twiddle_data[0][1][3]~q ),
	.twiddle_data014(\twiddle_data[0][1][4]~q ),
	.twiddle_data015(\twiddle_data[0][1][5]~q ),
	.twiddle_data016(\twiddle_data[0][1][6]~q ),
	.twiddle_data017(\twiddle_data[0][1][7]~q ),
	.twiddle_data007(\twiddle_data[0][0][7]~q ),
	.twiddle_data107(\twiddle_data[1][0][7]~q ),
	.twiddle_data110(\twiddle_data[1][1][0]~q ),
	.twiddle_data111(\twiddle_data[1][1][1]~q ),
	.twiddle_data112(\twiddle_data[1][1][2]~q ),
	.twiddle_data113(\twiddle_data[1][1][3]~q ),
	.twiddle_data114(\twiddle_data[1][1][4]~q ),
	.twiddle_data115(\twiddle_data[1][1][5]~q ),
	.twiddle_data116(\twiddle_data[1][1][6]~q ),
	.twiddle_data117(\twiddle_data[1][1][7]~q ),
	.twiddle_data207(\twiddle_data[2][0][7]~q ),
	.twiddle_data210(\twiddle_data[2][1][0]~q ),
	.twiddle_data211(\twiddle_data[2][1][1]~q ),
	.twiddle_data212(\twiddle_data[2][1][2]~q ),
	.twiddle_data213(\twiddle_data[2][1][3]~q ),
	.twiddle_data214(\twiddle_data[2][1][4]~q ),
	.twiddle_data215(\twiddle_data[2][1][5]~q ),
	.twiddle_data216(\twiddle_data[2][1][6]~q ),
	.twiddle_data217(\twiddle_data[2][1][7]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.slb_last_0(\gen_dft_1:bfpc|slb_last[0]~q ),
	.slb_last_1(\gen_dft_1:bfpc|slb_last[1]~q ),
	.slb_last_2(\gen_dft_1:bfpc|slb_last[2]~q ),
	.lut_out_tmp_0(\gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[0]~q ),
	.lut_out_tmp_1(\gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[1]~q ),
	.lut_out_tmp_2(\gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[2]~q ),
	.tdl_arr_3_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_4_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_5_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_6_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_2_1(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_11(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_12(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_13(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_14(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_15(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_1_1(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_11(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_12(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_13(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_14(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_15(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_0_1(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_11(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_12(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_13(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_14(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_15(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][0]~q ),
	.twiddle_data000(\twiddle_data[0][0][0]~q ),
	.twiddle_data001(\twiddle_data[0][0][1]~q ),
	.twiddle_data002(\twiddle_data[0][0][2]~q ),
	.twiddle_data003(\twiddle_data[0][0][3]~q ),
	.twiddle_data004(\twiddle_data[0][0][4]~q ),
	.twiddle_data005(\twiddle_data[0][0][5]~q ),
	.twiddle_data006(\twiddle_data[0][0][6]~q ),
	.twiddle_data100(\twiddle_data[1][0][0]~q ),
	.twiddle_data101(\twiddle_data[1][0][1]~q ),
	.twiddle_data102(\twiddle_data[1][0][2]~q ),
	.twiddle_data103(\twiddle_data[1][0][3]~q ),
	.twiddle_data104(\twiddle_data[1][0][4]~q ),
	.twiddle_data105(\twiddle_data[1][0][5]~q ),
	.twiddle_data106(\twiddle_data[1][0][6]~q ),
	.twiddle_data200(\twiddle_data[2][0][0]~q ),
	.twiddle_data201(\twiddle_data[2][0][1]~q ),
	.twiddle_data202(\twiddle_data[2][0][2]~q ),
	.twiddle_data203(\twiddle_data[2][0][3]~q ),
	.twiddle_data204(\twiddle_data[2][0][4]~q ),
	.twiddle_data205(\twiddle_data[2][0][5]~q ),
	.twiddle_data206(\twiddle_data[2][0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_bfp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_5_1(\ram_cxb_bfp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_2_1(\ram_cxb_bfp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_1(\ram_cxb_bfp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_1(\ram_cxb_bfp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_6_3(\ram_cxb_bfp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_5_3(\ram_cxb_bfp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_2_3(\ram_cxb_bfp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_bfp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_4_3(\ram_cxb_bfp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_6_0(\ram_cxb_bfp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_5_0(\ram_cxb_bfp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_2_0(\ram_cxb_bfp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\ram_cxb_bfp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_0(\ram_cxb_bfp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_6_2(\ram_cxb_bfp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_5_2(\ram_cxb_bfp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_2_2(\ram_cxb_bfp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_3_2(\ram_cxb_bfp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_4_2(\ram_cxb_bfp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_7_1(\ram_cxb_bfp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_bfp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_bfp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_bfp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_bfp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_6_5(\ram_cxb_bfp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_3_5(\ram_cxb_bfp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_4_5(\ram_cxb_bfp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_5_5(\ram_cxb_bfp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_7_7(\ram_cxb_bfp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_6_7(\ram_cxb_bfp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_3_7(\ram_cxb_bfp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_4_7(\ram_cxb_bfp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_5_7(\ram_cxb_bfp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_7_4(\ram_cxb_bfp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_6_4(\ram_cxb_bfp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_3_4(\ram_cxb_bfp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_4_4(\ram_cxb_bfp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_5_4(\ram_cxb_bfp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_7_6(\ram_cxb_bfp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_6_6(\ram_cxb_bfp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_3_6(\ram_cxb_bfp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_4_6(\ram_cxb_bfp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_5_6(\ram_cxb_bfp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_2_5(\ram_cxb_bfp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_bfp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_bfp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_bfp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_0_2(\ram_cxb_bfp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_1_2(\ram_cxb_bfp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_0_0(\ram_cxb_bfp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\ram_cxb_bfp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_0_7(\ram_cxb_bfp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_1_7(\ram_cxb_bfp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_5(\ram_cxb_bfp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_1_5(\ram_cxb_bfp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_bfp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_1_3(\ram_cxb_bfp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_1(\ram_cxb_bfp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_1(\ram_cxb_bfp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_bfp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_1_6(\ram_cxb_bfp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_4(\ram_cxb_bfp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_1_4(\ram_cxb_bfp_data|ram_in_reg[4][1]~q ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_cxb_data_r_1 ram_cxb_bfp_data(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_6_1(\ram_cxb_bfp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_5_1(\ram_cxb_bfp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_2_1(\ram_cxb_bfp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_1(\ram_cxb_bfp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_4_1(\ram_cxb_bfp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_6_3(\ram_cxb_bfp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_5_3(\ram_cxb_bfp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_2_3(\ram_cxb_bfp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_bfp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_4_3(\ram_cxb_bfp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_6_0(\ram_cxb_bfp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_5_0(\ram_cxb_bfp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_2_0(\ram_cxb_bfp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\ram_cxb_bfp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_4_0(\ram_cxb_bfp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_6_2(\ram_cxb_bfp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_5_2(\ram_cxb_bfp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_2_2(\ram_cxb_bfp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_3_2(\ram_cxb_bfp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_4_2(\ram_cxb_bfp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_7_1(\ram_cxb_bfp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_3(\ram_cxb_bfp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_bfp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_bfp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_bfp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_6_5(\ram_cxb_bfp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_3_5(\ram_cxb_bfp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_4_5(\ram_cxb_bfp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_5_5(\ram_cxb_bfp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_7_7(\ram_cxb_bfp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_6_7(\ram_cxb_bfp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_3_7(\ram_cxb_bfp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_4_7(\ram_cxb_bfp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_5_7(\ram_cxb_bfp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_7_4(\ram_cxb_bfp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_6_4(\ram_cxb_bfp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_3_4(\ram_cxb_bfp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_4_4(\ram_cxb_bfp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_5_4(\ram_cxb_bfp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_7_6(\ram_cxb_bfp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_6_6(\ram_cxb_bfp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_3_6(\ram_cxb_bfp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_4_6(\ram_cxb_bfp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_5_6(\ram_cxb_bfp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_2_5(\ram_cxb_bfp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_bfp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_bfp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_bfp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_0_2(\ram_cxb_bfp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_1_2(\ram_cxb_bfp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_0_0(\ram_cxb_bfp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\ram_cxb_bfp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_0_7(\ram_cxb_bfp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_1_7(\ram_cxb_bfp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_0_5(\ram_cxb_bfp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_1_5(\ram_cxb_bfp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_bfp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_1_3(\ram_cxb_bfp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_1(\ram_cxb_bfp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_1(\ram_cxb_bfp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_0_6(\ram_cxb_bfp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_1_6(\ram_cxb_bfp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_4(\ram_cxb_bfp_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_1_4(\ram_cxb_bfp_data|ram_in_reg[4][1]~q ),
	.ram_data_out1_14(\ccc|ram_data_out1[14]~q ),
	.ram_data_out2_14(\ccc|ram_data_out2[14]~q ),
	.ram_data_out3_14(\ccc|ram_data_out3[14]~q ),
	.ram_data_out0_14(\ccc|ram_data_out0[14]~q ),
	.sw_r_tdl_0_4(\sw_r_tdl[4][0]~q ),
	.sw_r_tdl_1_4(\sw_r_tdl[4][1]~q ),
	.ram_data_out1_13(\ccc|ram_data_out1[13]~q ),
	.ram_data_out2_13(\ccc|ram_data_out2[13]~q ),
	.ram_data_out3_13(\ccc|ram_data_out3[13]~q ),
	.ram_data_out0_13(\ccc|ram_data_out0[13]~q ),
	.ram_data_out1_10(\ccc|ram_data_out1[10]~q ),
	.ram_data_out2_10(\ccc|ram_data_out2[10]~q ),
	.ram_data_out3_10(\ccc|ram_data_out3[10]~q ),
	.ram_data_out0_10(\ccc|ram_data_out0[10]~q ),
	.ram_data_out1_11(\ccc|ram_data_out1[11]~q ),
	.ram_data_out2_11(\ccc|ram_data_out2[11]~q ),
	.ram_data_out3_11(\ccc|ram_data_out3[11]~q ),
	.ram_data_out0_11(\ccc|ram_data_out0[11]~q ),
	.ram_data_out1_12(\ccc|ram_data_out1[12]~q ),
	.ram_data_out2_12(\ccc|ram_data_out2[12]~q ),
	.ram_data_out3_12(\ccc|ram_data_out3[12]~q ),
	.ram_data_out0_12(\ccc|ram_data_out0[12]~q ),
	.ram_data_out1_15(\ccc|ram_data_out1[15]~q ),
	.ram_data_out2_15(\ccc|ram_data_out2[15]~q ),
	.ram_data_out3_15(\ccc|ram_data_out3[15]~q ),
	.ram_data_out0_15(\ccc|ram_data_out0[15]~q ),
	.ram_data_out1_7(\ccc|ram_data_out1[7]~q ),
	.ram_data_out2_7(\ccc|ram_data_out2[7]~q ),
	.ram_data_out3_7(\ccc|ram_data_out3[7]~q ),
	.ram_data_out0_7(\ccc|ram_data_out0[7]~q ),
	.ram_data_out1_6(\ccc|ram_data_out1[6]~q ),
	.ram_data_out2_6(\ccc|ram_data_out2[6]~q ),
	.ram_data_out3_6(\ccc|ram_data_out3[6]~q ),
	.ram_data_out0_6(\ccc|ram_data_out0[6]~q ),
	.ram_data_out1_3(\ccc|ram_data_out1[3]~q ),
	.ram_data_out2_3(\ccc|ram_data_out2[3]~q ),
	.ram_data_out3_3(\ccc|ram_data_out3[3]~q ),
	.ram_data_out0_3(\ccc|ram_data_out0[3]~q ),
	.ram_data_out1_4(\ccc|ram_data_out1[4]~q ),
	.ram_data_out2_4(\ccc|ram_data_out2[4]~q ),
	.ram_data_out3_4(\ccc|ram_data_out3[4]~q ),
	.ram_data_out0_4(\ccc|ram_data_out0[4]~q ),
	.ram_data_out1_5(\ccc|ram_data_out1[5]~q ),
	.ram_data_out2_5(\ccc|ram_data_out2[5]~q ),
	.ram_data_out3_5(\ccc|ram_data_out3[5]~q ),
	.ram_data_out0_5(\ccc|ram_data_out0[5]~q ),
	.ram_data_out1_2(\ccc|ram_data_out1[2]~q ),
	.ram_data_out2_2(\ccc|ram_data_out2[2]~q ),
	.ram_data_out3_2(\ccc|ram_data_out3[2]~q ),
	.ram_data_out0_2(\ccc|ram_data_out0[2]~q ),
	.ram_data_out2_8(\ccc|ram_data_out2[8]~q ),
	.ram_data_out3_8(\ccc|ram_data_out3[8]~q ),
	.ram_data_out0_8(\ccc|ram_data_out0[8]~q ),
	.ram_data_out1_8(\ccc|ram_data_out1[8]~q ),
	.ram_data_out2_9(\ccc|ram_data_out2[9]~q ),
	.ram_data_out3_9(\ccc|ram_data_out3[9]~q ),
	.ram_data_out0_9(\ccc|ram_data_out0[9]~q ),
	.ram_data_out1_9(\ccc|ram_data_out1[9]~q ),
	.ram_data_out3_0(\ccc|ram_data_out3[0]~q ),
	.ram_data_out0_0(\ccc|ram_data_out0[0]~q ),
	.ram_data_out1_0(\ccc|ram_data_out1[0]~q ),
	.ram_data_out2_0(\ccc|ram_data_out2[0]~q ),
	.ram_data_out3_1(\ccc|ram_data_out3[1]~q ),
	.ram_data_out0_1(\ccc|ram_data_out0[1]~q ),
	.ram_data_out1_1(\ccc|ram_data_out1[1]~q ),
	.ram_data_out2_1(\ccc|ram_data_out2[1]~q ),
	.clk(clk));

IFFT_asj_fft_cxb_data ram_cxb_wr_data(
	.reg_no_twiddle603(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][3]~q ),
	.reg_no_twiddle607(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][7]~q ),
	.reg_no_twiddle617(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][7]~q ),
	.reg_no_twiddle613(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][3]~q ),
	.reg_no_twiddle604(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][4]~q ),
	.reg_no_twiddle614(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][4]~q ),
	.reg_no_twiddle605(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][5]~q ),
	.reg_no_twiddle615(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][5]~q ),
	.reg_no_twiddle606(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][6]~q ),
	.reg_no_twiddle616(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][6]~q ),
	.reg_no_twiddle602(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][2]~q ),
	.ram_block6a3(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a3~portbdataout ),
	.ram_block6a2(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a2~portbdataout ),
	.reg_no_twiddle612(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][2]~q ),
	.reg_no_twiddle601(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][1]~q ),
	.reg_no_twiddle611(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][1]~q ),
	.reg_no_twiddle600(\gen_dft_1:bfpdft|reg_no_twiddle[6][0][0]~q ),
	.reg_no_twiddle610(\gen_dft_1:bfpdft|reg_no_twiddle[6][1][0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.tdl_arr_3_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][7]~q ),
	.tdl_arr_3_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][3]~q ),
	.tdl_arr_7_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][7]~q ),
	.tdl_arr_4_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][4]~q ),
	.tdl_arr_4_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][4]~q ),
	.tdl_arr_5_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][5]~q ),
	.tdl_arr_5_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][5]~q ),
	.tdl_arr_6_1(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_11(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_12(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_13(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_14(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][6]~q ),
	.tdl_arr_6_15(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][6]~q ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.tdl_arr_2_1(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_11(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_12(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_13(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_14(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][2]~q ),
	.tdl_arr_2_15(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][2]~q ),
	.ram_in_reg_1_3(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_2(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.tdl_arr_1_1(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_11(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_12(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_13(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_14(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][1]~q ),
	.tdl_arr_1_15(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_0(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.tdl_arr_0_1(\gen_dft_1:bfpdft|gen_da2:cm3|imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_11(\gen_dft_1:bfpdft|gen_da2:cm1|imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_12(\gen_dft_1:bfpdft|gen_da2:cm2|imag_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_13(\gen_dft_1:bfpdft|gen_da2:cm3|real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_14(\gen_dft_1:bfpdft|gen_da2:cm1|real_delay|tdl_arr[1][0]~q ),
	.tdl_arr_0_15(\gen_dft_1:bfpdft|gen_da2:cm2|real_delay|tdl_arr[1][0]~q ),
	.clk(clk));

IFFT_asj_fft_cxb_addr_1 \gen_wrsw_1:ram_cxb_wr (
	.ram_block6a0(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ),
	.ram_block6a1(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ),
	.ram_block6a01(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ),
	.ram_block6a11(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_3(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_0_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_2(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_0(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_0_01(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_11(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_31(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_11(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_21(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_01(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.clk(clk));

IFFT_asj_fft_wrswgen \gen_wrsw_1:get_wr_swtiches (
	.ram_block6a3(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a3~portbdataout ),
	.ram_block6a2(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a2~portbdataout ),
	.ram_block6a0(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ),
	.ram_block6a1(\gen_wrsw_1:get_wr_swtiches|swa_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.p_tdl_0_0(\p_tdl[0][0]~q ),
	.p_tdl_1_0(\p_tdl[0][1]~q ),
	.k_count_1(\gen_le256_mk:ctrl|k_count[1]~q ),
	.k_count_3(\gen_le256_mk:ctrl|k_count[3]~q ),
	.k_count_0(\gen_le256_mk:ctrl|k_count[0]~q ),
	.k_count_2(\gen_le256_mk:ctrl|k_count[2]~q ),
	.clk(clk));

IFFT_asj_fft_cxb_addr_2 ram_cxb_rd(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_2_0(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_0(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_0_0(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_1(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_3(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_1(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_2(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_0(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.rd_addr_d_2(\rd_adgen|rd_addr_d[2]~q ),
	.rd_addr_d_3(\rd_adgen|rd_addr_d[3]~q ),
	.rd_addr_d_0(\rd_adgen|rd_addr_d[0]~q ),
	.sw_0(\rd_adgen|sw[0]~q ),
	.rd_addr_c_0(\rd_adgen|rd_addr_c[0]~q ),
	.rd_addr_b_1(\rd_adgen|rd_addr_b[1]~q ),
	.sw_1(\rd_adgen|sw[1]~q ),
	.rd_addr_d_1(\rd_adgen|rd_addr_d[1]~q ),
	.clk(clk));

IFFT_asj_fft_dataadgen rd_adgen(
	.p_0(\gen_le256_mk:ctrl|p[0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.p_1(\gen_le256_mk:ctrl|p[1]~q ),
	.k_count_1(\gen_le256_mk:ctrl|k_count[1]~q ),
	.k_count_3(\gen_le256_mk:ctrl|k_count[3]~q ),
	.k_count_0(\gen_le256_mk:ctrl|k_count[0]~q ),
	.k_count_2(\gen_le256_mk:ctrl|k_count[2]~q ),
	.rd_addr_d_2(\rd_adgen|rd_addr_d[2]~q ),
	.rd_addr_d_3(\rd_adgen|rd_addr_d[3]~q ),
	.rd_addr_d_0(\rd_adgen|rd_addr_d[0]~q ),
	.sw_0(\rd_adgen|sw[0]~q ),
	.rd_addr_c_0(\rd_adgen|rd_addr_c[0]~q ),
	.rd_addr_b_1(\rd_adgen|rd_addr_b[1]~q ),
	.sw_1(\rd_adgen|sw[1]~q ),
	.rd_addr_d_1(\rd_adgen|rd_addr_d[1]~q ),
	.Mux1(\rd_adgen|Mux1~1_combout ),
	.Mux0(\rd_adgen|Mux0~1_combout ),
	.Mux11(\rd_adgen|Mux1~2_combout ),
	.Mux01(\rd_adgen|Mux0~2_combout ),
	.clk(clk));

IFFT_asj_fft_tdl_bit_rst_8 delay_ctrl_np(
	.next_pass_i(\gen_le256_mk:ctrl|next_pass_i~q ),
	.tdl_arr_9(\delay_ctrl_np|tdl_arr[9]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_m_k_counter \gen_le256_mk:ctrl (
	.blk_done_int1(\gen_le256_mk:ctrl|blk_done_int~q ),
	.next_block(\writer|next_block~q ),
	.p_0(\gen_le256_mk:ctrl|p[0]~q ),
	.data_rdy_vec_4(\data_rdy_vec[4]~q ),
	.next_pass_i1(\gen_le256_mk:ctrl|next_pass_i~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.p_1(\gen_le256_mk:ctrl|p[1]~q ),
	.k_count_1(\gen_le256_mk:ctrl|k_count[1]~q ),
	.k_count_3(\gen_le256_mk:ctrl|k_count[3]~q ),
	.k_count_0(\gen_le256_mk:ctrl|k_count[0]~q ),
	.k_count_2(\gen_le256_mk:ctrl|k_count[2]~q ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_auk_dspip_avalon_streaming_controller auk_dsp_interface_controller_1(
	.sink_in_work(\sink_in_work~q ),
	.at_source_valid_s(at_source_valid_s),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.sink_stall(\auk_dsp_atlantic_sink_1|sink_stall~combout ),
	.sink_stall_reg1(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.source_stall_reg1(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_ready_ctrl(\auk_dsp_interface_controller_1|sink_ready_ctrl~0_combout ),
	.master_sink_ena(\master_sink_ena~q ),
	.send_eop_s(\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.packet_error_s_1(\auk_dsp_atlantic_sink_1|packet_error_s[1]~q ),
	.packet_error_s_0(\auk_dsp_atlantic_sink_1|packet_error_s[0]~q ),
	.stall_controller_comb(\auk_dsp_atlantic_source_1|stall_controller_comb~0_combout ),
	.stall_reg1(\auk_dsp_interface_controller_1|stall_reg~q ),
	.sink_ready_ctrl1(\auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~0_combout ),
	.Mux01(\auk_dsp_atlantic_source_1|Mux0~1_combout ),
	.Mux02(\auk_dsp_atlantic_source_1|Mux0~2_combout ),
	.stall_controller_comb1(\auk_dsp_atlantic_source_1|stall_controller_comb~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_auk_dspip_avalon_streaming_source auk_dsp_atlantic_source_1(
	.at_source_data_14(at_source_data_14),
	.at_source_data_15(at_source_data_15),
	.at_source_data_16(at_source_data_16),
	.at_source_data_17(at_source_data_17),
	.at_source_data_18(at_source_data_18),
	.at_source_data_19(at_source_data_19),
	.at_source_data_20(at_source_data_20),
	.at_source_data_21(at_source_data_21),
	.at_source_data_6(at_source_data_6),
	.at_source_data_7(at_source_data_7),
	.at_source_data_8(at_source_data_8),
	.at_source_data_9(at_source_data_9),
	.at_source_data_10(at_source_data_10),
	.at_source_data_11(at_source_data_11),
	.at_source_data_12(at_source_data_12),
	.at_source_data_13(at_source_data_13),
	.at_source_data_0(at_source_data_0),
	.at_source_data_1(at_source_data_1),
	.at_source_data_2(at_source_data_2),
	.at_source_data_3(at_source_data_3),
	.at_source_data_4(at_source_data_4),
	.at_source_data_5(at_source_data_5),
	.master_source_ena(\master_source_ena~q ),
	.data({\fft_real_out[7]~q ,\fft_real_out[6]~q ,\fft_real_out[5]~q ,\fft_real_out[4]~q ,\fft_real_out[3]~q ,\fft_real_out[2]~q ,\fft_real_out[1]~q ,\fft_real_out[0]~q ,\fft_imag_out[7]~q ,\fft_imag_out[6]~q ,\fft_imag_out[5]~q ,\fft_imag_out[4]~q ,\fft_imag_out[3]~q ,
\fft_imag_out[2]~q ,\fft_imag_out[1]~q ,\fft_imag_out[0]~q ,\exponent_out[5]~q ,\exponent_out[4]~q ,\exponent_out[3]~q ,\exponent_out[2]~q ,\exponent_out[1]~q ,\exponent_out[0]~q }),
	.at_source_valid_s1(at_source_valid_s),
	.at_source_error_0(at_source_error_0),
	.at_source_error_1(at_source_error_1),
	.at_source_sop_s1(at_source_sop_s),
	.at_source_eop_s1(at_source_eop_s),
	.source_packet_error_1(\auk_dsp_interface_controller_1|source_packet_error[1]~q ),
	.source_packet_error_0(\auk_dsp_interface_controller_1|source_packet_error[0]~q ),
	.sink_stall_reg(\auk_dsp_interface_controller_1|sink_stall_reg~q ),
	.source_stall_reg(\auk_dsp_interface_controller_1|source_stall_reg~q ),
	.sink_ready_ctrl_d(\sink_ready_ctrl_d~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.sop(\sop~q ),
	.stall_controller_comb(\auk_dsp_atlantic_source_1|stall_controller_comb~0_combout ),
	.data_count({\data_count_sig[5]~q ,\data_count_sig[4]~q ,\data_count_sig[3]~q ,\data_count_sig[2]~q ,\data_count_sig[1]~q ,\data_count_sig[0]~q }),
	.source_stall_int_d1(\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.stall_reg(\auk_dsp_interface_controller_1|stall_reg~q ),
	.Mux0(\auk_dsp_atlantic_source_1|Mux0~0_combout ),
	.Mux01(\auk_dsp_atlantic_source_1|Mux0~1_combout ),
	.Mux02(\auk_dsp_atlantic_source_1|Mux0~2_combout ),
	.stall_controller_comb1(\auk_dsp_atlantic_source_1|stall_controller_comb~1_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready));

IFFT_asj_fft_4dp_ram_2 dat_A(
	.q_b_14(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_141(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_13(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_131(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_10(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_11(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_12(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_15(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_151(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_7(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_6(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_3(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_4(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_5(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_2(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_8(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_9(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_0(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_1(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_16(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_17(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_18(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.wren_a_1(\wren_a[1]~q ),
	.a_ram_data_in_bus_46(\ccc|a_ram_data_in_bus[46]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_9(\ccc|wraddress_a_bus[9]~q ),
	.wraddress_a_bus_10(\ccc|wraddress_a_bus[10]~q ),
	.wraddress_a_bus_11(\ccc|wraddress_a_bus[11]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_9(\ccc|rdaddress_a_bus[9]~q ),
	.rdaddress_a_bus_10(\ccc|rdaddress_a_bus[10]~q ),
	.rdaddress_a_bus_11(\ccc|rdaddress_a_bus[11]~q ),
	.wren_a_2(\wren_a[2]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.wraddress_a_bus_12(\ccc|wraddress_a_bus[12]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.rdaddress_a_bus_12(\ccc|rdaddress_a_bus[12]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.wren_a_3(\wren_a[3]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.wren_a_0(\wren_a[0]~q ),
	.a_ram_data_in_bus_62(\ccc|a_ram_data_in_bus[62]~q ),
	.wraddress_a_bus_13(\ccc|wraddress_a_bus[13]~q ),
	.rdaddress_a_bus_13(\ccc|rdaddress_a_bus[13]~q ),
	.a_ram_data_in_bus_45(\ccc|a_ram_data_in_bus[45]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_61(\ccc|a_ram_data_in_bus[61]~q ),
	.a_ram_data_in_bus_42(\ccc|a_ram_data_in_bus[42]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.a_ram_data_in_bus_58(\ccc|a_ram_data_in_bus[58]~q ),
	.a_ram_data_in_bus_43(\ccc|a_ram_data_in_bus[43]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_59(\ccc|a_ram_data_in_bus[59]~q ),
	.a_ram_data_in_bus_44(\ccc|a_ram_data_in_bus[44]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.a_ram_data_in_bus_60(\ccc|a_ram_data_in_bus[60]~q ),
	.a_ram_data_in_bus_47(\ccc|a_ram_data_in_bus[47]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_63(\ccc|a_ram_data_in_bus[63]~q ),
	.a_ram_data_in_bus_39(\ccc|a_ram_data_in_bus[39]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_55(\ccc|a_ram_data_in_bus[55]~q ),
	.a_ram_data_in_bus_38(\ccc|a_ram_data_in_bus[38]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_54(\ccc|a_ram_data_in_bus[54]~q ),
	.a_ram_data_in_bus_35(\ccc|a_ram_data_in_bus[35]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_51(\ccc|a_ram_data_in_bus[51]~q ),
	.a_ram_data_in_bus_36(\ccc|a_ram_data_in_bus[36]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_52(\ccc|a_ram_data_in_bus[52]~q ),
	.a_ram_data_in_bus_37(\ccc|a_ram_data_in_bus[37]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_53(\ccc|a_ram_data_in_bus[53]~q ),
	.a_ram_data_in_bus_34(\ccc|a_ram_data_in_bus[34]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_50(\ccc|a_ram_data_in_bus[50]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_56(\ccc|a_ram_data_in_bus[56]~q ),
	.a_ram_data_in_bus_40(\ccc|a_ram_data_in_bus[40]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_57(\ccc|a_ram_data_in_bus[57]~q ),
	.a_ram_data_in_bus_41(\ccc|a_ram_data_in_bus[41]~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.a_ram_data_in_bus_48(\ccc|a_ram_data_in_bus[48]~q ),
	.a_ram_data_in_bus_32(\ccc|a_ram_data_in_bus[32]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_49(\ccc|a_ram_data_in_bus[49]~q ),
	.a_ram_data_in_bus_33(\ccc|a_ram_data_in_bus[33]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk));

IFFT_asj_fft_cnt_ctrl ccc(
	.ram_block6a0(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ),
	.ram_block6a1(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ),
	.data_rdy_vec_10(\data_rdy_vec[10]~q ),
	.q_b_14(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_141(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_144(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_145(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_146(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_147(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_13(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_131(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_134(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_135(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_136(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_137(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_10(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_104(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_105(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_106(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_107(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_11(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_114(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_115(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_116(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_117(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_12(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_124(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_125(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_126(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_127(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_15(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_151(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_154(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_155(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_156(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_157(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_7(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_74(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_75(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_76(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_77(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_6(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_64(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_65(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_66(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_67(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_3(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_34(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_35(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_36(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_37(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_4(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_44(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_45(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_46(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_47(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_5(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_54(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_55(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_56(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_57(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_2(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_24(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_25(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_26(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_27(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_8(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_84(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_85(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_86(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_87(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_9(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_94(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_95(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_96(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_97(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_0(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_04(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_05(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_06(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_07(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_1(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_16(\dat_A|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_17(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_18(\dat_A|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_19(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_110(\dat_A|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_118(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_119(\dat_A|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.b_ram_data_in_bus_46(\ccc|b_ram_data_in_bus[46]~q ),
	.wraddress_b_bus_0(\ccc|wraddress_b_bus[0]~q ),
	.wraddress_b_bus_9(\ccc|wraddress_b_bus[9]~q ),
	.wraddress_b_bus_10(\ccc|wraddress_b_bus[10]~q ),
	.wraddress_b_bus_11(\ccc|wraddress_b_bus[11]~q ),
	.rdaddress_b_bus_0(\ccc|rdaddress_b_bus[0]~q ),
	.rdaddress_b_bus_9(\ccc|rdaddress_b_bus[9]~q ),
	.rdaddress_b_bus_10(\ccc|rdaddress_b_bus[10]~q ),
	.rdaddress_b_bus_11(\ccc|rdaddress_b_bus[11]~q ),
	.a_ram_data_in_bus_46(\ccc|a_ram_data_in_bus[46]~q ),
	.wraddress_a_bus_0(\ccc|wraddress_a_bus[0]~q ),
	.wraddress_a_bus_9(\ccc|wraddress_a_bus[9]~q ),
	.wraddress_a_bus_10(\ccc|wraddress_a_bus[10]~q ),
	.wraddress_a_bus_11(\ccc|wraddress_a_bus[11]~q ),
	.rdaddress_a_bus_0(\ccc|rdaddress_a_bus[0]~q ),
	.rdaddress_a_bus_9(\ccc|rdaddress_a_bus[9]~q ),
	.rdaddress_a_bus_10(\ccc|rdaddress_a_bus[10]~q ),
	.rdaddress_a_bus_11(\ccc|rdaddress_a_bus[11]~q ),
	.b_ram_data_in_bus_30(\ccc|b_ram_data_in_bus[30]~q ),
	.wraddress_b_bus_12(\ccc|wraddress_b_bus[12]~q ),
	.wraddress_b_bus_5(\ccc|wraddress_b_bus[5]~q ),
	.rdaddress_b_bus_12(\ccc|rdaddress_b_bus[12]~q ),
	.rdaddress_b_bus_5(\ccc|rdaddress_b_bus[5]~q ),
	.a_ram_data_in_bus_30(\ccc|a_ram_data_in_bus[30]~q ),
	.wraddress_a_bus_12(\ccc|wraddress_a_bus[12]~q ),
	.wraddress_a_bus_5(\ccc|wraddress_a_bus[5]~q ),
	.rdaddress_a_bus_12(\ccc|rdaddress_a_bus[12]~q ),
	.rdaddress_a_bus_5(\ccc|rdaddress_a_bus[5]~q ),
	.b_ram_data_in_bus_14(\ccc|b_ram_data_in_bus[14]~q ),
	.wraddress_b_bus_1(\ccc|wraddress_b_bus[1]~q ),
	.rdaddress_b_bus_1(\ccc|rdaddress_b_bus[1]~q ),
	.a_ram_data_in_bus_14(\ccc|a_ram_data_in_bus[14]~q ),
	.wraddress_a_bus_1(\ccc|wraddress_a_bus[1]~q ),
	.rdaddress_a_bus_1(\ccc|rdaddress_a_bus[1]~q ),
	.b_ram_data_in_bus_62(\ccc|b_ram_data_in_bus[62]~q ),
	.wraddress_b_bus_13(\ccc|wraddress_b_bus[13]~q ),
	.rdaddress_b_bus_13(\ccc|rdaddress_b_bus[13]~q ),
	.a_ram_data_in_bus_62(\ccc|a_ram_data_in_bus[62]~q ),
	.wraddress_a_bus_13(\ccc|wraddress_a_bus[13]~q ),
	.rdaddress_a_bus_13(\ccc|rdaddress_a_bus[13]~q ),
	.b_ram_data_in_bus_45(\ccc|b_ram_data_in_bus[45]~q ),
	.a_ram_data_in_bus_45(\ccc|a_ram_data_in_bus[45]~q ),
	.b_ram_data_in_bus_29(\ccc|b_ram_data_in_bus[29]~q ),
	.a_ram_data_in_bus_29(\ccc|a_ram_data_in_bus[29]~q ),
	.b_ram_data_in_bus_13(\ccc|b_ram_data_in_bus[13]~q ),
	.a_ram_data_in_bus_13(\ccc|a_ram_data_in_bus[13]~q ),
	.b_ram_data_in_bus_61(\ccc|b_ram_data_in_bus[61]~q ),
	.a_ram_data_in_bus_61(\ccc|a_ram_data_in_bus[61]~q ),
	.b_ram_data_in_bus_42(\ccc|b_ram_data_in_bus[42]~q ),
	.a_ram_data_in_bus_42(\ccc|a_ram_data_in_bus[42]~q ),
	.b_ram_data_in_bus_26(\ccc|b_ram_data_in_bus[26]~q ),
	.a_ram_data_in_bus_26(\ccc|a_ram_data_in_bus[26]~q ),
	.b_ram_data_in_bus_10(\ccc|b_ram_data_in_bus[10]~q ),
	.a_ram_data_in_bus_10(\ccc|a_ram_data_in_bus[10]~q ),
	.b_ram_data_in_bus_58(\ccc|b_ram_data_in_bus[58]~q ),
	.a_ram_data_in_bus_58(\ccc|a_ram_data_in_bus[58]~q ),
	.b_ram_data_in_bus_43(\ccc|b_ram_data_in_bus[43]~q ),
	.a_ram_data_in_bus_43(\ccc|a_ram_data_in_bus[43]~q ),
	.b_ram_data_in_bus_27(\ccc|b_ram_data_in_bus[27]~q ),
	.a_ram_data_in_bus_27(\ccc|a_ram_data_in_bus[27]~q ),
	.b_ram_data_in_bus_11(\ccc|b_ram_data_in_bus[11]~q ),
	.a_ram_data_in_bus_11(\ccc|a_ram_data_in_bus[11]~q ),
	.b_ram_data_in_bus_59(\ccc|b_ram_data_in_bus[59]~q ),
	.a_ram_data_in_bus_59(\ccc|a_ram_data_in_bus[59]~q ),
	.b_ram_data_in_bus_44(\ccc|b_ram_data_in_bus[44]~q ),
	.a_ram_data_in_bus_44(\ccc|a_ram_data_in_bus[44]~q ),
	.b_ram_data_in_bus_28(\ccc|b_ram_data_in_bus[28]~q ),
	.a_ram_data_in_bus_28(\ccc|a_ram_data_in_bus[28]~q ),
	.b_ram_data_in_bus_12(\ccc|b_ram_data_in_bus[12]~q ),
	.a_ram_data_in_bus_12(\ccc|a_ram_data_in_bus[12]~q ),
	.b_ram_data_in_bus_60(\ccc|b_ram_data_in_bus[60]~q ),
	.a_ram_data_in_bus_60(\ccc|a_ram_data_in_bus[60]~q ),
	.b_ram_data_in_bus_47(\ccc|b_ram_data_in_bus[47]~q ),
	.a_ram_data_in_bus_47(\ccc|a_ram_data_in_bus[47]~q ),
	.b_ram_data_in_bus_31(\ccc|b_ram_data_in_bus[31]~q ),
	.a_ram_data_in_bus_31(\ccc|a_ram_data_in_bus[31]~q ),
	.b_ram_data_in_bus_15(\ccc|b_ram_data_in_bus[15]~q ),
	.a_ram_data_in_bus_15(\ccc|a_ram_data_in_bus[15]~q ),
	.b_ram_data_in_bus_63(\ccc|b_ram_data_in_bus[63]~q ),
	.a_ram_data_in_bus_63(\ccc|a_ram_data_in_bus[63]~q ),
	.b_ram_data_in_bus_39(\ccc|b_ram_data_in_bus[39]~q ),
	.a_ram_data_in_bus_39(\ccc|a_ram_data_in_bus[39]~q ),
	.b_ram_data_in_bus_23(\ccc|b_ram_data_in_bus[23]~q ),
	.a_ram_data_in_bus_23(\ccc|a_ram_data_in_bus[23]~q ),
	.b_ram_data_in_bus_7(\ccc|b_ram_data_in_bus[7]~q ),
	.a_ram_data_in_bus_7(\ccc|a_ram_data_in_bus[7]~q ),
	.b_ram_data_in_bus_55(\ccc|b_ram_data_in_bus[55]~q ),
	.a_ram_data_in_bus_55(\ccc|a_ram_data_in_bus[55]~q ),
	.b_ram_data_in_bus_38(\ccc|b_ram_data_in_bus[38]~q ),
	.a_ram_data_in_bus_38(\ccc|a_ram_data_in_bus[38]~q ),
	.b_ram_data_in_bus_22(\ccc|b_ram_data_in_bus[22]~q ),
	.a_ram_data_in_bus_22(\ccc|a_ram_data_in_bus[22]~q ),
	.b_ram_data_in_bus_6(\ccc|b_ram_data_in_bus[6]~q ),
	.a_ram_data_in_bus_6(\ccc|a_ram_data_in_bus[6]~q ),
	.b_ram_data_in_bus_54(\ccc|b_ram_data_in_bus[54]~q ),
	.a_ram_data_in_bus_54(\ccc|a_ram_data_in_bus[54]~q ),
	.b_ram_data_in_bus_35(\ccc|b_ram_data_in_bus[35]~q ),
	.a_ram_data_in_bus_35(\ccc|a_ram_data_in_bus[35]~q ),
	.b_ram_data_in_bus_19(\ccc|b_ram_data_in_bus[19]~q ),
	.a_ram_data_in_bus_19(\ccc|a_ram_data_in_bus[19]~q ),
	.b_ram_data_in_bus_3(\ccc|b_ram_data_in_bus[3]~q ),
	.a_ram_data_in_bus_3(\ccc|a_ram_data_in_bus[3]~q ),
	.b_ram_data_in_bus_51(\ccc|b_ram_data_in_bus[51]~q ),
	.a_ram_data_in_bus_51(\ccc|a_ram_data_in_bus[51]~q ),
	.b_ram_data_in_bus_36(\ccc|b_ram_data_in_bus[36]~q ),
	.a_ram_data_in_bus_36(\ccc|a_ram_data_in_bus[36]~q ),
	.b_ram_data_in_bus_20(\ccc|b_ram_data_in_bus[20]~q ),
	.a_ram_data_in_bus_20(\ccc|a_ram_data_in_bus[20]~q ),
	.b_ram_data_in_bus_4(\ccc|b_ram_data_in_bus[4]~q ),
	.a_ram_data_in_bus_4(\ccc|a_ram_data_in_bus[4]~q ),
	.b_ram_data_in_bus_52(\ccc|b_ram_data_in_bus[52]~q ),
	.a_ram_data_in_bus_52(\ccc|a_ram_data_in_bus[52]~q ),
	.b_ram_data_in_bus_37(\ccc|b_ram_data_in_bus[37]~q ),
	.a_ram_data_in_bus_37(\ccc|a_ram_data_in_bus[37]~q ),
	.b_ram_data_in_bus_21(\ccc|b_ram_data_in_bus[21]~q ),
	.a_ram_data_in_bus_21(\ccc|a_ram_data_in_bus[21]~q ),
	.b_ram_data_in_bus_5(\ccc|b_ram_data_in_bus[5]~q ),
	.a_ram_data_in_bus_5(\ccc|a_ram_data_in_bus[5]~q ),
	.b_ram_data_in_bus_53(\ccc|b_ram_data_in_bus[53]~q ),
	.a_ram_data_in_bus_53(\ccc|a_ram_data_in_bus[53]~q ),
	.b_ram_data_in_bus_34(\ccc|b_ram_data_in_bus[34]~q ),
	.a_ram_data_in_bus_34(\ccc|a_ram_data_in_bus[34]~q ),
	.b_ram_data_in_bus_18(\ccc|b_ram_data_in_bus[18]~q ),
	.a_ram_data_in_bus_18(\ccc|a_ram_data_in_bus[18]~q ),
	.b_ram_data_in_bus_2(\ccc|b_ram_data_in_bus[2]~q ),
	.a_ram_data_in_bus_2(\ccc|a_ram_data_in_bus[2]~q ),
	.b_ram_data_in_bus_50(\ccc|b_ram_data_in_bus[50]~q ),
	.a_ram_data_in_bus_50(\ccc|a_ram_data_in_bus[50]~q ),
	.b_ram_data_in_bus_24(\ccc|b_ram_data_in_bus[24]~q ),
	.a_ram_data_in_bus_24(\ccc|a_ram_data_in_bus[24]~q ),
	.b_ram_data_in_bus_8(\ccc|b_ram_data_in_bus[8]~q ),
	.a_ram_data_in_bus_8(\ccc|a_ram_data_in_bus[8]~q ),
	.b_ram_data_in_bus_56(\ccc|b_ram_data_in_bus[56]~q ),
	.a_ram_data_in_bus_56(\ccc|a_ram_data_in_bus[56]~q ),
	.b_ram_data_in_bus_40(\ccc|b_ram_data_in_bus[40]~q ),
	.a_ram_data_in_bus_40(\ccc|a_ram_data_in_bus[40]~q ),
	.b_ram_data_in_bus_25(\ccc|b_ram_data_in_bus[25]~q ),
	.a_ram_data_in_bus_25(\ccc|a_ram_data_in_bus[25]~q ),
	.b_ram_data_in_bus_9(\ccc|b_ram_data_in_bus[9]~q ),
	.a_ram_data_in_bus_9(\ccc|a_ram_data_in_bus[9]~q ),
	.b_ram_data_in_bus_57(\ccc|b_ram_data_in_bus[57]~q ),
	.a_ram_data_in_bus_57(\ccc|a_ram_data_in_bus[57]~q ),
	.b_ram_data_in_bus_41(\ccc|b_ram_data_in_bus[41]~q ),
	.a_ram_data_in_bus_41(\ccc|a_ram_data_in_bus[41]~q ),
	.b_ram_data_in_bus_0(\ccc|b_ram_data_in_bus[0]~q ),
	.a_ram_data_in_bus_0(\ccc|a_ram_data_in_bus[0]~q ),
	.b_ram_data_in_bus_48(\ccc|b_ram_data_in_bus[48]~q ),
	.a_ram_data_in_bus_48(\ccc|a_ram_data_in_bus[48]~q ),
	.b_ram_data_in_bus_32(\ccc|b_ram_data_in_bus[32]~q ),
	.a_ram_data_in_bus_32(\ccc|a_ram_data_in_bus[32]~q ),
	.b_ram_data_in_bus_16(\ccc|b_ram_data_in_bus[16]~q ),
	.a_ram_data_in_bus_16(\ccc|a_ram_data_in_bus[16]~q ),
	.b_ram_data_in_bus_1(\ccc|b_ram_data_in_bus[1]~q ),
	.a_ram_data_in_bus_1(\ccc|a_ram_data_in_bus[1]~q ),
	.b_ram_data_in_bus_49(\ccc|b_ram_data_in_bus[49]~q ),
	.a_ram_data_in_bus_49(\ccc|a_ram_data_in_bus[49]~q ),
	.b_ram_data_in_bus_33(\ccc|b_ram_data_in_bus[33]~q ),
	.a_ram_data_in_bus_33(\ccc|a_ram_data_in_bus[33]~q ),
	.b_ram_data_in_bus_17(\ccc|b_ram_data_in_bus[17]~q ),
	.a_ram_data_in_bus_17(\ccc|a_ram_data_in_bus[17]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_0_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_3(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_0_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_1_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_1_2(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_2_01(\ram_cxb_rd|ram_in_reg[0][2]~q ),
	.ram_in_reg_3_01(\ram_cxb_rd|ram_in_reg[0][3]~q ),
	.ram_in_reg_1_31(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_01(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_11(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_21(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_01(\ram_cxb_rd|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_11(\ram_cxb_rd|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_32(\ram_cxb_rd|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_12(\ram_cxb_rd|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_22(\ram_cxb_rd|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_02(\ram_cxb_rd|ram_in_reg[0][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_02(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_12(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.ram_data_out1_14(\ccc|ram_data_out1[14]~q ),
	.ram_data_out2_14(\ccc|ram_data_out2[14]~q ),
	.ram_data_out3_14(\ccc|ram_data_out3[14]~q ),
	.ram_data_out0_14(\ccc|ram_data_out0[14]~q ),
	.ram_data_out1_13(\ccc|ram_data_out1[13]~q ),
	.ram_data_out2_13(\ccc|ram_data_out2[13]~q ),
	.ram_data_out3_13(\ccc|ram_data_out3[13]~q ),
	.ram_data_out0_13(\ccc|ram_data_out0[13]~q ),
	.ram_data_out1_10(\ccc|ram_data_out1[10]~q ),
	.ram_data_out2_10(\ccc|ram_data_out2[10]~q ),
	.ram_data_out3_10(\ccc|ram_data_out3[10]~q ),
	.ram_data_out0_10(\ccc|ram_data_out0[10]~q ),
	.ram_data_out1_11(\ccc|ram_data_out1[11]~q ),
	.ram_data_out2_11(\ccc|ram_data_out2[11]~q ),
	.ram_data_out3_11(\ccc|ram_data_out3[11]~q ),
	.ram_data_out0_11(\ccc|ram_data_out0[11]~q ),
	.ram_data_out1_12(\ccc|ram_data_out1[12]~q ),
	.ram_data_out2_12(\ccc|ram_data_out2[12]~q ),
	.ram_data_out3_12(\ccc|ram_data_out3[12]~q ),
	.ram_data_out0_12(\ccc|ram_data_out0[12]~q ),
	.ram_data_out1_15(\ccc|ram_data_out1[15]~q ),
	.ram_data_out2_15(\ccc|ram_data_out2[15]~q ),
	.ram_data_out3_15(\ccc|ram_data_out3[15]~q ),
	.ram_data_out0_15(\ccc|ram_data_out0[15]~q ),
	.ram_data_out1_7(\ccc|ram_data_out1[7]~q ),
	.ram_data_out2_7(\ccc|ram_data_out2[7]~q ),
	.ram_data_out3_7(\ccc|ram_data_out3[7]~q ),
	.ram_data_out0_7(\ccc|ram_data_out0[7]~q ),
	.ram_data_out1_6(\ccc|ram_data_out1[6]~q ),
	.ram_data_out2_6(\ccc|ram_data_out2[6]~q ),
	.ram_data_out3_6(\ccc|ram_data_out3[6]~q ),
	.ram_data_out0_6(\ccc|ram_data_out0[6]~q ),
	.ram_data_out1_3(\ccc|ram_data_out1[3]~q ),
	.ram_data_out2_3(\ccc|ram_data_out2[3]~q ),
	.ram_data_out3_3(\ccc|ram_data_out3[3]~q ),
	.ram_data_out0_3(\ccc|ram_data_out0[3]~q ),
	.ram_data_out1_4(\ccc|ram_data_out1[4]~q ),
	.ram_data_out2_4(\ccc|ram_data_out2[4]~q ),
	.ram_data_out3_4(\ccc|ram_data_out3[4]~q ),
	.ram_data_out0_4(\ccc|ram_data_out0[4]~q ),
	.ram_data_out1_5(\ccc|ram_data_out1[5]~q ),
	.ram_data_out2_5(\ccc|ram_data_out2[5]~q ),
	.ram_data_out3_5(\ccc|ram_data_out3[5]~q ),
	.ram_data_out0_5(\ccc|ram_data_out0[5]~q ),
	.ram_data_out1_2(\ccc|ram_data_out1[2]~q ),
	.ram_data_out2_2(\ccc|ram_data_out2[2]~q ),
	.ram_data_out3_2(\ccc|ram_data_out3[2]~q ),
	.ram_data_out0_2(\ccc|ram_data_out0[2]~q ),
	.ram_data_out2_8(\ccc|ram_data_out2[8]~q ),
	.ram_data_out3_8(\ccc|ram_data_out3[8]~q ),
	.ram_data_out0_8(\ccc|ram_data_out0[8]~q ),
	.ram_data_out1_8(\ccc|ram_data_out1[8]~q ),
	.ram_data_out2_9(\ccc|ram_data_out2[9]~q ),
	.ram_data_out3_9(\ccc|ram_data_out3[9]~q ),
	.ram_data_out0_9(\ccc|ram_data_out0[9]~q ),
	.ram_data_out1_9(\ccc|ram_data_out1[9]~q ),
	.ram_data_out3_0(\ccc|ram_data_out3[0]~q ),
	.ram_data_out0_0(\ccc|ram_data_out0[0]~q ),
	.ram_data_out1_0(\ccc|ram_data_out1[0]~q ),
	.ram_data_out2_0(\ccc|ram_data_out2[0]~q ),
	.ram_data_out3_1(\ccc|ram_data_out3[1]~q ),
	.ram_data_out0_1(\ccc|ram_data_out0[1]~q ),
	.ram_data_out1_1(\ccc|ram_data_out1[1]~q ),
	.ram_data_out2_1(\ccc|ram_data_out2[1]~q ),
	.ram_a_not_b_vec_10(\ram_a_not_b_vec[10]~q ),
	.ram_a_not_b_vec_1(\ram_a_not_b_vec[1]~q ),
	.sel_anb_addr(\sel_anb_addr~combout ),
	.clk(clk));

IFFT_asj_fft_in_write_sgl writer(
	.next_block1(\writer|next_block~q ),
	.data_rdy_int1(\writer|data_rdy_int~q ),
	.wren_1(\writer|wren[1]~q ),
	.data_in_r_6(\writer|data_in_r[6]~q ),
	.wr_address_i_int_0(\writer|wr_address_i_int[0]~q ),
	.wr_address_i_int_1(\writer|wr_address_i_int[1]~q ),
	.wr_address_i_int_2(\writer|wr_address_i_int[2]~q ),
	.wr_address_i_int_3(\writer|wr_address_i_int[3]~q ),
	.wren_2(\writer|wren[2]~q ),
	.wren_3(\writer|wren[3]~q ),
	.wren_0(\writer|wren[0]~q ),
	.data_in_r_5(\writer|data_in_r[5]~q ),
	.data_in_r_2(\writer|data_in_r[2]~q ),
	.data_in_r_3(\writer|data_in_r[3]~q ),
	.data_in_r_4(\writer|data_in_r[4]~q ),
	.data_in_r_7(\writer|data_in_r[7]~q ),
	.data_in_i_7(\writer|data_in_i[7]~q ),
	.data_in_i_6(\writer|data_in_i[6]~q ),
	.data_in_i_3(\writer|data_in_i[3]~q ),
	.data_in_i_4(\writer|data_in_i[4]~q ),
	.data_in_i_5(\writer|data_in_i[5]~q ),
	.data_in_i_2(\writer|data_in_i[2]~q ),
	.data_in_r_0(\writer|data_in_r[0]~q ),
	.data_in_r_1(\writer|data_in_r[1]~q ),
	.data_in_i_0(\writer|data_in_i[0]~q ),
	.data_in_i_1(\writer|data_in_i[1]~q ),
	.core_real_in_6(\core_real_in[6]~q ),
	.core_real_in_5(\core_real_in[5]~q ),
	.core_real_in_2(\core_real_in[2]~q ),
	.core_real_in_3(\core_real_in[3]~q ),
	.core_real_in_4(\core_real_in[4]~q ),
	.core_real_in_7(\core_real_in[7]~q ),
	.core_imag_in_7(\core_imag_in[7]~q ),
	.core_imag_in_6(\core_imag_in[6]~q ),
	.core_imag_in_3(\core_imag_in[3]~q ),
	.core_imag_in_4(\core_imag_in[4]~q ),
	.core_imag_in_5(\core_imag_in[5]~q ),
	.core_imag_in_2(\core_imag_in[2]~q ),
	.core_real_in_0(\core_real_in[0]~q ),
	.core_real_in_1(\core_real_in[1]~q ),
	.core_imag_in_0(\core_imag_in[0]~q ),
	.core_imag_in_1(\core_imag_in[1]~q ),
	.anb1(\writer|anb~q ),
	.send_sop_s(\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_wrengen sel_we(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.wc_i1(\sel_we|wc_i~q ),
	.wd_i1(\sel_we|wd_i~q ),
	.ram_a_not_b_vec_26(\ram_a_not_b_vec[26]~q ),
	.p_cd_en_0(\p_cd_en[0]~q ),
	.p_cd_en_1(\p_cd_en[1]~q ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_4dp_ram_3 dat_B(
	.q_b_14(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_141(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_13(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_131(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_10(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_11(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_12(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_15(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_151(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_7(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_6(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_3(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_4(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_5(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_2(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_8(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_9(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_0(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_1(\dat_B|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_16(\dat_B|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_17(\dat_B|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_18(\dat_B|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.wren_b_1(\wren_b[1]~q ),
	.b_ram_data_in_bus_46(\ccc|b_ram_data_in_bus[46]~q ),
	.wraddress_b_bus_0(\ccc|wraddress_b_bus[0]~q ),
	.wraddress_b_bus_9(\ccc|wraddress_b_bus[9]~q ),
	.wraddress_b_bus_10(\ccc|wraddress_b_bus[10]~q ),
	.wraddress_b_bus_11(\ccc|wraddress_b_bus[11]~q ),
	.rdaddress_b_bus_0(\ccc|rdaddress_b_bus[0]~q ),
	.rdaddress_b_bus_9(\ccc|rdaddress_b_bus[9]~q ),
	.rdaddress_b_bus_10(\ccc|rdaddress_b_bus[10]~q ),
	.rdaddress_b_bus_11(\ccc|rdaddress_b_bus[11]~q ),
	.wren_b_2(\wren_b[2]~q ),
	.b_ram_data_in_bus_30(\ccc|b_ram_data_in_bus[30]~q ),
	.wraddress_b_bus_12(\ccc|wraddress_b_bus[12]~q ),
	.wraddress_b_bus_5(\ccc|wraddress_b_bus[5]~q ),
	.rdaddress_b_bus_12(\ccc|rdaddress_b_bus[12]~q ),
	.rdaddress_b_bus_5(\ccc|rdaddress_b_bus[5]~q ),
	.wren_b_3(\wren_b[3]~q ),
	.b_ram_data_in_bus_14(\ccc|b_ram_data_in_bus[14]~q ),
	.wraddress_b_bus_1(\ccc|wraddress_b_bus[1]~q ),
	.rdaddress_b_bus_1(\ccc|rdaddress_b_bus[1]~q ),
	.wren_b_0(\wren_b[0]~q ),
	.b_ram_data_in_bus_62(\ccc|b_ram_data_in_bus[62]~q ),
	.wraddress_b_bus_13(\ccc|wraddress_b_bus[13]~q ),
	.rdaddress_b_bus_13(\ccc|rdaddress_b_bus[13]~q ),
	.b_ram_data_in_bus_45(\ccc|b_ram_data_in_bus[45]~q ),
	.b_ram_data_in_bus_29(\ccc|b_ram_data_in_bus[29]~q ),
	.b_ram_data_in_bus_13(\ccc|b_ram_data_in_bus[13]~q ),
	.b_ram_data_in_bus_61(\ccc|b_ram_data_in_bus[61]~q ),
	.b_ram_data_in_bus_42(\ccc|b_ram_data_in_bus[42]~q ),
	.b_ram_data_in_bus_26(\ccc|b_ram_data_in_bus[26]~q ),
	.b_ram_data_in_bus_10(\ccc|b_ram_data_in_bus[10]~q ),
	.b_ram_data_in_bus_58(\ccc|b_ram_data_in_bus[58]~q ),
	.b_ram_data_in_bus_43(\ccc|b_ram_data_in_bus[43]~q ),
	.b_ram_data_in_bus_27(\ccc|b_ram_data_in_bus[27]~q ),
	.b_ram_data_in_bus_11(\ccc|b_ram_data_in_bus[11]~q ),
	.b_ram_data_in_bus_59(\ccc|b_ram_data_in_bus[59]~q ),
	.b_ram_data_in_bus_44(\ccc|b_ram_data_in_bus[44]~q ),
	.b_ram_data_in_bus_28(\ccc|b_ram_data_in_bus[28]~q ),
	.b_ram_data_in_bus_12(\ccc|b_ram_data_in_bus[12]~q ),
	.b_ram_data_in_bus_60(\ccc|b_ram_data_in_bus[60]~q ),
	.b_ram_data_in_bus_47(\ccc|b_ram_data_in_bus[47]~q ),
	.b_ram_data_in_bus_31(\ccc|b_ram_data_in_bus[31]~q ),
	.b_ram_data_in_bus_15(\ccc|b_ram_data_in_bus[15]~q ),
	.b_ram_data_in_bus_63(\ccc|b_ram_data_in_bus[63]~q ),
	.b_ram_data_in_bus_39(\ccc|b_ram_data_in_bus[39]~q ),
	.b_ram_data_in_bus_23(\ccc|b_ram_data_in_bus[23]~q ),
	.b_ram_data_in_bus_7(\ccc|b_ram_data_in_bus[7]~q ),
	.b_ram_data_in_bus_55(\ccc|b_ram_data_in_bus[55]~q ),
	.b_ram_data_in_bus_38(\ccc|b_ram_data_in_bus[38]~q ),
	.b_ram_data_in_bus_22(\ccc|b_ram_data_in_bus[22]~q ),
	.b_ram_data_in_bus_6(\ccc|b_ram_data_in_bus[6]~q ),
	.b_ram_data_in_bus_54(\ccc|b_ram_data_in_bus[54]~q ),
	.b_ram_data_in_bus_35(\ccc|b_ram_data_in_bus[35]~q ),
	.b_ram_data_in_bus_19(\ccc|b_ram_data_in_bus[19]~q ),
	.b_ram_data_in_bus_3(\ccc|b_ram_data_in_bus[3]~q ),
	.b_ram_data_in_bus_51(\ccc|b_ram_data_in_bus[51]~q ),
	.b_ram_data_in_bus_36(\ccc|b_ram_data_in_bus[36]~q ),
	.b_ram_data_in_bus_20(\ccc|b_ram_data_in_bus[20]~q ),
	.b_ram_data_in_bus_4(\ccc|b_ram_data_in_bus[4]~q ),
	.b_ram_data_in_bus_52(\ccc|b_ram_data_in_bus[52]~q ),
	.b_ram_data_in_bus_37(\ccc|b_ram_data_in_bus[37]~q ),
	.b_ram_data_in_bus_21(\ccc|b_ram_data_in_bus[21]~q ),
	.b_ram_data_in_bus_5(\ccc|b_ram_data_in_bus[5]~q ),
	.b_ram_data_in_bus_53(\ccc|b_ram_data_in_bus[53]~q ),
	.b_ram_data_in_bus_34(\ccc|b_ram_data_in_bus[34]~q ),
	.b_ram_data_in_bus_18(\ccc|b_ram_data_in_bus[18]~q ),
	.b_ram_data_in_bus_2(\ccc|b_ram_data_in_bus[2]~q ),
	.b_ram_data_in_bus_50(\ccc|b_ram_data_in_bus[50]~q ),
	.b_ram_data_in_bus_24(\ccc|b_ram_data_in_bus[24]~q ),
	.b_ram_data_in_bus_8(\ccc|b_ram_data_in_bus[8]~q ),
	.b_ram_data_in_bus_56(\ccc|b_ram_data_in_bus[56]~q ),
	.b_ram_data_in_bus_40(\ccc|b_ram_data_in_bus[40]~q ),
	.b_ram_data_in_bus_25(\ccc|b_ram_data_in_bus[25]~q ),
	.b_ram_data_in_bus_9(\ccc|b_ram_data_in_bus[9]~q ),
	.b_ram_data_in_bus_57(\ccc|b_ram_data_in_bus[57]~q ),
	.b_ram_data_in_bus_41(\ccc|b_ram_data_in_bus[41]~q ),
	.b_ram_data_in_bus_0(\ccc|b_ram_data_in_bus[0]~q ),
	.b_ram_data_in_bus_48(\ccc|b_ram_data_in_bus[48]~q ),
	.b_ram_data_in_bus_32(\ccc|b_ram_data_in_bus[32]~q ),
	.b_ram_data_in_bus_16(\ccc|b_ram_data_in_bus[16]~q ),
	.b_ram_data_in_bus_1(\ccc|b_ram_data_in_bus[1]~q ),
	.b_ram_data_in_bus_49(\ccc|b_ram_data_in_bus[49]~q ),
	.b_ram_data_in_bus_33(\ccc|b_ram_data_in_bus[33]~q ),
	.b_ram_data_in_bus_17(\ccc|b_ram_data_in_bus[17]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk));

IFFT_asj_fft_4dp_ram \gen_M4K_Output:dat_C (
	.q_b_10(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_2(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_11(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_3(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_12(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_4(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_13(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_131(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_5(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_14(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_141(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_6(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_15(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_151(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_7(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.wc_vec_3(\wc_vec[3]~q ),
	.ram_block6a0(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ),
	.ram_block6a1(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ),
	.rdaddress_c_bus_0(\rdaddress_c_bus[0]~q ),
	.rdaddress_c_bus_13(\rdaddress_c_bus[13]~q ),
	.rdaddress_c_bus_10(\rdaddress_c_bus[10]~q ),
	.rdaddress_c_bus_3(\rdaddress_c_bus[3]~q ),
	.rdaddress_c_bus_14(\rdaddress_c_bus[14]~q ),
	.rdaddress_c_bus_15(\rdaddress_c_bus[15]~q ),
	.rdaddress_c_bus_11(\rdaddress_c_bus[11]~q ),
	.rdaddress_c_bus_7(\rdaddress_c_bus[7]~q ),
	.q_b_9(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_1(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_16(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_17(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_18(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_8(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_0(\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_0_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_3(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_0_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_1_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_1_2(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_1_31(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_01(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_11(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_21(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_01(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_11(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.clk(clk));

IFFT_asj_fft_4dp_ram_1 \gen_M4K_Output:dat_D (
	.q_b_10(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_101(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_102(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_103(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_2(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_21(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_22(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_23(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_11(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_111(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_112(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_113(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_3(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_31(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_32(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_33(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_12(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_121(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_122(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_123(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_4(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_41(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_42(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_43(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_13(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_131(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_132(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_133(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_5(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_51(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_52(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_53(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_14(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_141(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_142(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_143(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_6(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_61(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_62(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_63(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_15(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_151(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_152(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_153(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_7(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_71(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_72(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.q_b_73(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.ram_block6a0(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0~portbdataout ),
	.ram_block6a1(\gen_wrsw_1:ram_cxb_wr|sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1~portbdataout ),
	.rdaddress_c_bus_0(\rdaddress_c_bus[0]~q ),
	.rdaddress_c_bus_13(\rdaddress_c_bus[13]~q ),
	.rdaddress_c_bus_10(\rdaddress_c_bus[10]~q ),
	.rdaddress_c_bus_3(\rdaddress_c_bus[3]~q ),
	.wd_vec_3(\wd_vec[3]~q ),
	.rdaddress_c_bus_14(\rdaddress_c_bus[14]~q ),
	.rdaddress_c_bus_15(\rdaddress_c_bus[15]~q ),
	.rdaddress_c_bus_11(\rdaddress_c_bus[11]~q ),
	.rdaddress_c_bus_7(\rdaddress_c_bus[7]~q ),
	.q_b_9(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_91(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_92(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_93(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_1(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_16(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_17(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_18(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_8(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_81(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_82(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_83(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_0(\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_01(\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_02(\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_03(\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_2_3(\ram_cxb_wr_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_0_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][0]~q ),
	.ram_in_reg_1_3(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[3][1]~q ),
	.ram_in_reg_2_0(\ram_cxb_wr_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_0_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_1(\ram_cxb_wr_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_1_1(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[1][1]~q ),
	.ram_in_reg_2_2(\ram_cxb_wr_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_1_2(\gen_wrsw_1:ram_cxb_wr|ram_in_reg[2][1]~q ),
	.ram_in_reg_2_7(\ram_cxb_wr_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_4(\ram_cxb_wr_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_2_5(\ram_cxb_wr_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_6(\ram_cxb_wr_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_3_3(\ram_cxb_wr_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_0(\ram_cxb_wr_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_1(\ram_cxb_wr_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_2(\ram_cxb_wr_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_7(\ram_cxb_wr_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_4(\ram_cxb_wr_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_3_5(\ram_cxb_wr_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_6(\ram_cxb_wr_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_4_3(\ram_cxb_wr_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_0(\ram_cxb_wr_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_1(\ram_cxb_wr_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_2(\ram_cxb_wr_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_7(\ram_cxb_wr_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_4(\ram_cxb_wr_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_4_5(\ram_cxb_wr_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_6(\ram_cxb_wr_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_5_3(\ram_cxb_wr_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_0(\ram_cxb_wr_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_1(\ram_cxb_wr_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_2(\ram_cxb_wr_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_7(\ram_cxb_wr_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_4(\ram_cxb_wr_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_5_5(\ram_cxb_wr_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_6(\ram_cxb_wr_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_6_3(\ram_cxb_wr_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_0(\ram_cxb_wr_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_1(\ram_cxb_wr_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_2(\ram_cxb_wr_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_7(\ram_cxb_wr_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_4(\ram_cxb_wr_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_6_5(\ram_cxb_wr_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_6(\ram_cxb_wr_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_7_3(\ram_cxb_wr_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_0(\ram_cxb_wr_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_1(\ram_cxb_wr_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_2(\ram_cxb_wr_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_7(\ram_cxb_wr_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_4(\ram_cxb_wr_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_7_5(\ram_cxb_wr_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_6(\ram_cxb_wr_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_1_31(\ram_cxb_wr_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_01(\ram_cxb_wr_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_11(\ram_cxb_wr_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_21(\ram_cxb_wr_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_7(\ram_cxb_wr_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_4(\ram_cxb_wr_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_1_5(\ram_cxb_wr_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_6(\ram_cxb_wr_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_0_3(\ram_cxb_wr_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_01(\ram_cxb_wr_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_11(\ram_cxb_wr_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_2(\ram_cxb_wr_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_7(\ram_cxb_wr_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_4(\ram_cxb_wr_data|ram_in_reg[4][0]~q ),
	.ram_in_reg_0_5(\ram_cxb_wr_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_6(\ram_cxb_wr_data|ram_in_reg[6][0]~q ),
	.clk(clk));

IFFT_asj_fft_tdl_bit_rst_9 delay_lpp_en(
	.tdl_arr_5(\delay_lpp_en|tdl_arr[5]~q ),
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_lpp_serial \gen_radix_4_last_pass:lpp (
	.data_real_o_0(\gen_radix_4_last_pass:lpp|data_real_o[0]~q ),
	.data_real_o_1(\gen_radix_4_last_pass:lpp|data_real_o[1]~q ),
	.data_real_o_2(\gen_radix_4_last_pass:lpp|data_real_o[2]~q ),
	.data_real_o_3(\gen_radix_4_last_pass:lpp|data_real_o[3]~q ),
	.data_real_o_4(\gen_radix_4_last_pass:lpp|data_real_o[4]~q ),
	.data_real_o_5(\gen_radix_4_last_pass:lpp|data_real_o[5]~q ),
	.data_real_o_6(\gen_radix_4_last_pass:lpp|data_real_o[6]~q ),
	.data_real_o_7(\gen_radix_4_last_pass:lpp|data_real_o[7]~q ),
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.data_imag_o_0(\gen_radix_4_last_pass:lpp|data_imag_o[0]~q ),
	.data_imag_o_1(\gen_radix_4_last_pass:lpp|data_imag_o[1]~q ),
	.data_imag_o_2(\gen_radix_4_last_pass:lpp|data_imag_o[2]~q ),
	.data_imag_o_3(\gen_radix_4_last_pass:lpp|data_imag_o[3]~q ),
	.data_imag_o_4(\gen_radix_4_last_pass:lpp|data_imag_o[4]~q ),
	.data_imag_o_5(\gen_radix_4_last_pass:lpp|data_imag_o[5]~q ),
	.data_imag_o_6(\gen_radix_4_last_pass:lpp|data_imag_o[6]~q ),
	.data_imag_o_7(\gen_radix_4_last_pass:lpp|data_imag_o[7]~q ),
	.ram_in_reg_2_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][2]~q ),
	.data_3_real_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][6]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][4]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][2]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][0]~q }),
	.data_1_real_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][6]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][4]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][2]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][0]~q }),
	.data_3_imag_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][6]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][4]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][2]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][0]~q }),
	.data_1_imag_i({\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][7]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][6]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][5]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][4]~q ,
\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][3]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][2]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][1]~q ,\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][0]~q }),
	.ram_in_reg_3_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_4_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_5_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_6_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_7_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_1_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_0_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][0]~q ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_cxb_data_r \gen_radix_4_last_pass:ram_cxb_lpp_data (
	.lpp_ram_data_out_10_3(\lpp_ram_data_out[3][10]~q ),
	.lpp_ram_data_out_10_0(\lpp_ram_data_out[0][10]~q ),
	.lpp_ram_data_out_10_1(\lpp_ram_data_out[1][10]~q ),
	.lpp_ram_data_out_10_2(\lpp_ram_data_out[2][10]~q ),
	.tdl_arr_0_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.tdl_arr_1_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.lpp_ram_data_out_2_3(\lpp_ram_data_out[3][2]~q ),
	.lpp_ram_data_out_2_0(\lpp_ram_data_out[0][2]~q ),
	.lpp_ram_data_out_2_1(\lpp_ram_data_out[1][2]~q ),
	.lpp_ram_data_out_2_2(\lpp_ram_data_out[2][2]~q ),
	.lpp_ram_data_out_11_3(\lpp_ram_data_out[3][11]~q ),
	.lpp_ram_data_out_11_0(\lpp_ram_data_out[0][11]~q ),
	.lpp_ram_data_out_11_1(\lpp_ram_data_out[1][11]~q ),
	.lpp_ram_data_out_11_2(\lpp_ram_data_out[2][11]~q ),
	.lpp_ram_data_out_3_3(\lpp_ram_data_out[3][3]~q ),
	.lpp_ram_data_out_3_0(\lpp_ram_data_out[0][3]~q ),
	.lpp_ram_data_out_3_1(\lpp_ram_data_out[1][3]~q ),
	.lpp_ram_data_out_3_2(\lpp_ram_data_out[2][3]~q ),
	.lpp_ram_data_out_12_3(\lpp_ram_data_out[3][12]~q ),
	.lpp_ram_data_out_12_0(\lpp_ram_data_out[0][12]~q ),
	.lpp_ram_data_out_12_1(\lpp_ram_data_out[1][12]~q ),
	.lpp_ram_data_out_12_2(\lpp_ram_data_out[2][12]~q ),
	.lpp_ram_data_out_4_3(\lpp_ram_data_out[3][4]~q ),
	.lpp_ram_data_out_4_0(\lpp_ram_data_out[0][4]~q ),
	.lpp_ram_data_out_4_1(\lpp_ram_data_out[1][4]~q ),
	.lpp_ram_data_out_4_2(\lpp_ram_data_out[2][4]~q ),
	.lpp_ram_data_out_13_3(\lpp_ram_data_out[3][13]~q ),
	.lpp_ram_data_out_13_0(\lpp_ram_data_out[0][13]~q ),
	.lpp_ram_data_out_13_1(\lpp_ram_data_out[1][13]~q ),
	.lpp_ram_data_out_13_2(\lpp_ram_data_out[2][13]~q ),
	.lpp_ram_data_out_5_3(\lpp_ram_data_out[3][5]~q ),
	.lpp_ram_data_out_5_0(\lpp_ram_data_out[0][5]~q ),
	.lpp_ram_data_out_5_1(\lpp_ram_data_out[1][5]~q ),
	.lpp_ram_data_out_5_2(\lpp_ram_data_out[2][5]~q ),
	.lpp_ram_data_out_14_3(\lpp_ram_data_out[3][14]~q ),
	.lpp_ram_data_out_14_0(\lpp_ram_data_out[0][14]~q ),
	.lpp_ram_data_out_14_1(\lpp_ram_data_out[1][14]~q ),
	.lpp_ram_data_out_14_2(\lpp_ram_data_out[2][14]~q ),
	.lpp_ram_data_out_6_3(\lpp_ram_data_out[3][6]~q ),
	.lpp_ram_data_out_6_0(\lpp_ram_data_out[0][6]~q ),
	.lpp_ram_data_out_6_1(\lpp_ram_data_out[1][6]~q ),
	.lpp_ram_data_out_6_2(\lpp_ram_data_out[2][6]~q ),
	.lpp_ram_data_out_15_3(\lpp_ram_data_out[3][15]~q ),
	.lpp_ram_data_out_15_0(\lpp_ram_data_out[0][15]~q ),
	.lpp_ram_data_out_15_1(\lpp_ram_data_out[1][15]~q ),
	.lpp_ram_data_out_15_2(\lpp_ram_data_out[2][15]~q ),
	.lpp_ram_data_out_7_3(\lpp_ram_data_out[3][7]~q ),
	.lpp_ram_data_out_7_0(\lpp_ram_data_out[0][7]~q ),
	.lpp_ram_data_out_7_1(\lpp_ram_data_out[1][7]~q ),
	.lpp_ram_data_out_7_2(\lpp_ram_data_out[2][7]~q ),
	.lpp_ram_data_out_9_3(\lpp_ram_data_out[3][9]~q ),
	.lpp_ram_data_out_9_0(\lpp_ram_data_out[0][9]~q ),
	.lpp_ram_data_out_9_1(\lpp_ram_data_out[1][9]~q ),
	.lpp_ram_data_out_9_2(\lpp_ram_data_out[2][9]~q ),
	.lpp_ram_data_out_1_3(\lpp_ram_data_out[3][1]~q ),
	.lpp_ram_data_out_1_0(\lpp_ram_data_out[0][1]~q ),
	.lpp_ram_data_out_1_1(\lpp_ram_data_out[1][1]~q ),
	.lpp_ram_data_out_1_2(\lpp_ram_data_out[2][1]~q ),
	.lpp_ram_data_out_8_3(\lpp_ram_data_out[3][8]~q ),
	.lpp_ram_data_out_8_0(\lpp_ram_data_out[0][8]~q ),
	.lpp_ram_data_out_8_1(\lpp_ram_data_out[1][8]~q ),
	.lpp_ram_data_out_8_2(\lpp_ram_data_out[2][8]~q ),
	.lpp_ram_data_out_0_3(\lpp_ram_data_out[3][0]~q ),
	.lpp_ram_data_out_0_0(\lpp_ram_data_out[0][0]~q ),
	.lpp_ram_data_out_0_1(\lpp_ram_data_out[1][0]~q ),
	.lpp_ram_data_out_0_2(\lpp_ram_data_out[2][0]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_2_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][2]~q ),
	.ram_in_reg_2_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][2]~q ),
	.ram_in_reg_2_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][2]~q ),
	.ram_in_reg_2_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][2]~q ),
	.ram_in_reg_2_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][2]~q ),
	.ram_in_reg_2_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][2]~q ),
	.ram_in_reg_2_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][2]~q ),
	.ram_in_reg_2_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][2]~q ),
	.ram_in_reg_3_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][3]~q ),
	.ram_in_reg_3_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][3]~q ),
	.ram_in_reg_3_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][3]~q ),
	.ram_in_reg_3_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][3]~q ),
	.ram_in_reg_3_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][3]~q ),
	.ram_in_reg_3_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][3]~q ),
	.ram_in_reg_3_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][3]~q ),
	.ram_in_reg_4_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][4]~q ),
	.ram_in_reg_4_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][4]~q ),
	.ram_in_reg_4_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][4]~q ),
	.ram_in_reg_4_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][4]~q ),
	.ram_in_reg_4_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][4]~q ),
	.ram_in_reg_4_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][4]~q ),
	.ram_in_reg_4_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][4]~q ),
	.ram_in_reg_4_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][4]~q ),
	.ram_in_reg_5_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][5]~q ),
	.ram_in_reg_5_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][5]~q ),
	.ram_in_reg_5_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][5]~q ),
	.ram_in_reg_5_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][5]~q ),
	.ram_in_reg_5_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][5]~q ),
	.ram_in_reg_5_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][5]~q ),
	.ram_in_reg_5_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][5]~q ),
	.ram_in_reg_5_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][5]~q ),
	.ram_in_reg_6_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][6]~q ),
	.ram_in_reg_6_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][6]~q ),
	.ram_in_reg_6_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][6]~q ),
	.ram_in_reg_6_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][6]~q ),
	.ram_in_reg_6_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][6]~q ),
	.ram_in_reg_6_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][6]~q ),
	.ram_in_reg_6_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][6]~q ),
	.ram_in_reg_6_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][6]~q ),
	.ram_in_reg_7_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][7]~q ),
	.ram_in_reg_7_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][7]~q ),
	.ram_in_reg_7_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][7]~q ),
	.ram_in_reg_7_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][7]~q ),
	.ram_in_reg_7_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][7]~q ),
	.ram_in_reg_7_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][7]~q ),
	.ram_in_reg_7_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][7]~q ),
	.ram_in_reg_7_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][7]~q ),
	.ram_in_reg_1_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][1]~q ),
	.ram_in_reg_1_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][1]~q ),
	.ram_in_reg_1_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][1]~q ),
	.ram_in_reg_1_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][1]~q ),
	.ram_in_reg_1_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][1]~q ),
	.ram_in_reg_1_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][1]~q ),
	.ram_in_reg_1_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][1]~q ),
	.ram_in_reg_1_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][1]~q ),
	.ram_in_reg_0_3(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[3][0]~q ),
	.ram_in_reg_0_7(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[7][0]~q ),
	.ram_in_reg_0_1(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[1][0]~q ),
	.ram_in_reg_0_5(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[5][0]~q ),
	.ram_in_reg_0_2(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[2][0]~q ),
	.ram_in_reg_0_0(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[0][0]~q ),
	.ram_in_reg_0_6(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[6][0]~q ),
	.ram_in_reg_0_4(\gen_radix_4_last_pass:ram_cxb_lpp_data|ram_in_reg[4][0]~q ),
	.clk(clk));

IFFT_asj_fft_lpprdadgen \gen_radix_4_last_pass:gen_lpp_addr (
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.tdl_arr_19(\gen_dft_1:delay_blk_done2|tdl_arr[19]~q ),
	.data_rdy_int(\writer|data_rdy_int~q ),
	.tdl_arr_0_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][0]~q ),
	.tdl_arr_1_4(\gen_radix_4_last_pass:gen_lpp_addr|gen_M4K:delay_swd|tdl_arr[4][1]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.rd_addr_d_0(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[0]~q ),
	.rd_addr_d_1(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[1]~q ),
	.sw_0(\gen_radix_4_last_pass:gen_lpp_addr|sw[0]~q ),
	.sw_1(\gen_radix_4_last_pass:gen_lpp_addr|sw[1]~q ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_cxb_addr \gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp (
	.global_clock_enable(\global_clock_enable~0_combout ),
	.ram_in_reg_0_0(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ),
	.ram_in_reg_1_0(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ),
	.ram_in_reg_2_1(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[1][2]~q ),
	.ram_in_reg_3_3(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[3][3]~q ),
	.ram_in_reg_3_0(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ),
	.rd_addr_d_0(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[0]~q ),
	.rd_addr_d_1(\gen_radix_4_last_pass:gen_lpp_addr|rd_addr_d[1]~q ),
	.sw_0(\gen_radix_4_last_pass:gen_lpp_addr|sw[0]~q ),
	.sw_1(\gen_radix_4_last_pass:gen_lpp_addr|sw[1]~q ),
	.ram_in_reg_3_01(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][3]~_wirecell_combout ),
	.ram_in_reg_2_11(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[1][2]~_wirecell_combout ),
	.ram_in_reg_3_31(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[3][3]~_wirecell_combout ),
	.clk(clk));

IFFT_asj_fft_3dp_rom twrom(
	.q_a_0(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_1(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_2(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_3(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_4(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_5(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_6(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_7(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_01(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_11(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_21(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_31(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_41(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_51(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_61(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_71(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_02(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_12(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_22(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_32(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_42(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_52(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_62(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_72(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_03(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_13(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_23(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_33(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_43(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_53(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_63(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_73(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_04(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_14(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_24(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_34(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_44(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_54(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_64(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_74(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_a_05(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_a_15(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_a_25(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_a_35(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_a_45(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_a_55(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_a_65(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_a_75(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.twad_tdl_0_6(\twid_factors|twad_tdl[6][0]~q ),
	.twad_tdl_1_6(\twid_factors|twad_tdl[6][1]~q ),
	.twad_tdl_2_6(\twid_factors|twad_tdl[6][2]~q ),
	.twad_tdl_3_6(\twid_factors|twad_tdl[6][3]~q ),
	.clk(clk));

IFFT_asj_fft_twadgen twid_factors(
	.global_clock_enable(\global_clock_enable~0_combout ),
	.twad_tdl_0_6(\twid_factors|twad_tdl[6][0]~q ),
	.twad_tdl_1_6(\twid_factors|twad_tdl[6][1]~q ),
	.twad_tdl_2_6(\twid_factors|twad_tdl[6][2]~q ),
	.twad_tdl_3_6(\twid_factors|twad_tdl[6][3]~q ),
	.Mux1(\rd_adgen|Mux1~1_combout ),
	.Mux0(\rd_adgen|Mux0~1_combout ),
	.Mux11(\rd_adgen|Mux1~2_combout ),
	.Mux01(\rd_adgen|Mux0~2_combout ),
	.clk(clk));

IFFT_asj_fft_tdl_bit_rst_6 \gen_dft_1:delay_blk_done2 (
	.tdl_arr_11(\gen_dft_1:delay_blk_done|tdl_arr[11]~q ),
	.tdl_arr_19(\gen_dft_1:delay_blk_done2|tdl_arr[19]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_bfp_ctrl \gen_dft_1:bfpc (
	.tdl_arr_4(\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.tdl_arr_11(\gen_dft_1:delay_blk_done|tdl_arr[11]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.blk_exp_0(\gen_dft_1:bfpc|blk_exp[0]~q ),
	.blk_exp_1(\gen_dft_1:bfpc|blk_exp[1]~q ),
	.blk_exp_2(\gen_dft_1:bfpc|blk_exp[2]~q ),
	.blk_exp_3(\gen_dft_1:bfpc|blk_exp[3]~q ),
	.blk_exp_4(\gen_dft_1:bfpc|blk_exp[4]~q ),
	.blk_exp_5(\gen_dft_1:bfpc|blk_exp[5]~q ),
	.slb_last_0(\gen_dft_1:bfpc|slb_last[0]~q ),
	.slb_last_1(\gen_dft_1:bfpc|slb_last[1]~q ),
	.slb_last_2(\gen_dft_1:bfpc|slb_last[2]~q ),
	.lut_out_tmp_0(\gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[0]~q ),
	.lut_out_tmp_1(\gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[1]~q ),
	.lut_out_tmp_2(\gen_dft_1:bfpdft|gen_disc:bfp_detect|lut_out_tmp[2]~q ),
	.en_slb(\en_slb~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_tdl_bit_rst_5 \gen_dft_1:delay_blk_done (
	.blk_done_int(\gen_le256_mk:ctrl|blk_done_int~q ),
	.tdl_arr_11(\gen_dft_1:delay_blk_done|tdl_arr[11]~q ),
	.global_clock_enable(\global_clock_enable~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

dffeas sink_in_work(
	.clk(clk),
	.d(\sink_in_work~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_in_work~q ),
	.prn(vcc));
defparam sink_in_work.is_wysiwyg = "true";
defparam sink_in_work.power_up = "low";

dffeas master_source_ena(
	.clk(clk),
	.d(\oe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\master_source_ena~q ),
	.prn(vcc));
defparam master_source_ena.is_wysiwyg = "true";
defparam master_source_ena.power_up = "low";

dffeas \fft_real_out[0] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[0]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[0]~q ),
	.prn(vcc));
defparam \fft_real_out[0] .is_wysiwyg = "true";
defparam \fft_real_out[0] .power_up = "low";

dffeas \fft_real_out[1] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[1]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[1]~q ),
	.prn(vcc));
defparam \fft_real_out[1] .is_wysiwyg = "true";
defparam \fft_real_out[1] .power_up = "low";

dffeas \fft_real_out[2] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[2]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[2]~q ),
	.prn(vcc));
defparam \fft_real_out[2] .is_wysiwyg = "true";
defparam \fft_real_out[2] .power_up = "low";

dffeas \fft_real_out[3] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[3]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[3]~q ),
	.prn(vcc));
defparam \fft_real_out[3] .is_wysiwyg = "true";
defparam \fft_real_out[3] .power_up = "low";

dffeas \fft_real_out[4] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[4]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[4]~q ),
	.prn(vcc));
defparam \fft_real_out[4] .is_wysiwyg = "true";
defparam \fft_real_out[4] .power_up = "low";

dffeas \fft_real_out[5] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[5]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[5]~q ),
	.prn(vcc));
defparam \fft_real_out[5] .is_wysiwyg = "true";
defparam \fft_real_out[5] .power_up = "low";

dffeas \fft_real_out[6] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[6]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[6]~q ),
	.prn(vcc));
defparam \fft_real_out[6] .is_wysiwyg = "true";
defparam \fft_real_out[6] .power_up = "low";

dffeas \fft_real_out[7] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_real_o[7]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_imag_o[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_real_out[7]~q ),
	.prn(vcc));
defparam \fft_real_out[7] .is_wysiwyg = "true";
defparam \fft_real_out[7] .power_up = "low";

dffeas \fft_imag_out[0] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[0]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[0]~q ),
	.prn(vcc));
defparam \fft_imag_out[0] .is_wysiwyg = "true";
defparam \fft_imag_out[0] .power_up = "low";

dffeas \fft_imag_out[1] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[1]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[1]~q ),
	.prn(vcc));
defparam \fft_imag_out[1] .is_wysiwyg = "true";
defparam \fft_imag_out[1] .power_up = "low";

dffeas \fft_imag_out[2] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[2]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[2]~q ),
	.prn(vcc));
defparam \fft_imag_out[2] .is_wysiwyg = "true";
defparam \fft_imag_out[2] .power_up = "low";

dffeas \fft_imag_out[3] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[3]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[3]~q ),
	.prn(vcc));
defparam \fft_imag_out[3] .is_wysiwyg = "true";
defparam \fft_imag_out[3] .power_up = "low";

dffeas \fft_imag_out[4] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[4]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[4]~q ),
	.prn(vcc));
defparam \fft_imag_out[4] .is_wysiwyg = "true";
defparam \fft_imag_out[4] .power_up = "low";

dffeas \fft_imag_out[5] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[5]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[5]~q ),
	.prn(vcc));
defparam \fft_imag_out[5] .is_wysiwyg = "true";
defparam \fft_imag_out[5] .power_up = "low";

dffeas \fft_imag_out[6] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[6]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[6]~q ),
	.prn(vcc));
defparam \fft_imag_out[6] .is_wysiwyg = "true";
defparam \fft_imag_out[6] .power_up = "low";

dffeas \fft_imag_out[7] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:lpp|data_imag_o[7]~q ),
	.asdata(\gen_radix_4_last_pass:lpp|data_real_o[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\fft_imag_out[1]~0_combout ),
	.sload(\fft_dirn_stream~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_imag_out[7]~q ),
	.prn(vcc));
defparam \fft_imag_out[7] .is_wysiwyg = "true";
defparam \fft_imag_out[7] .power_up = "low";

dffeas oe(
	.clk(clk),
	.d(\WideNor1~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\oe~q ),
	.prn(vcc));
defparam oe.is_wysiwyg = "true";
defparam oe.power_up = "low";

dffeas fft_dirn_stream(
	.clk(clk),
	.d(\fft_dirn_stream~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_dirn_stream~q ),
	.prn(vcc));
defparam fft_dirn_stream.is_wysiwyg = "true";
defparam fft_dirn_stream.power_up = "low";

dffeas \fft_s2_cur.WAIT_FOR_LPP_INPUT (
	.clk(clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.prn(vcc));
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .is_wysiwyg = "true";
defparam \fft_s2_cur.WAIT_FOR_LPP_INPUT .power_up = "low";

dffeas sop_out(
	.clk(clk),
	.d(\fft_s2_cur.FIRST_LPP_C~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sop_out~q ),
	.prn(vcc));
defparam sop_out.is_wysiwyg = "true";
defparam sop_out.power_up = "low";

dffeas fft_dirn_held_o2(
	.clk(clk),
	.d(\fft_dirn_held_o2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_dirn_held_o2~q ),
	.prn(vcc));
defparam fft_dirn_held_o2.is_wysiwyg = "true";
defparam fft_dirn_held_o2.power_up = "low";

dffeas \lpp_count_offset[5] (
	.clk(clk),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~0_combout ),
	.q(\lpp_count_offset[5]~q ),
	.prn(vcc));
defparam \lpp_count_offset[5] .is_wysiwyg = "true";
defparam \lpp_count_offset[5] .power_up = "low";

dffeas \lpp_count_offset[1] (
	.clk(clk),
	.d(\Add1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~0_combout ),
	.q(\lpp_count_offset[1]~q ),
	.prn(vcc));
defparam \lpp_count_offset[1] .is_wysiwyg = "true";
defparam \lpp_count_offset[1] .power_up = "low";

dffeas \lpp_count_offset[2] (
	.clk(clk),
	.d(\Add1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~0_combout ),
	.q(\lpp_count_offset[2]~q ),
	.prn(vcc));
defparam \lpp_count_offset[2] .is_wysiwyg = "true";
defparam \lpp_count_offset[2] .power_up = "low";

dffeas \lpp_count_offset[3] (
	.clk(clk),
	.d(\Add1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~0_combout ),
	.q(\lpp_count_offset[3]~q ),
	.prn(vcc));
defparam \lpp_count_offset[3] .is_wysiwyg = "true";
defparam \lpp_count_offset[3] .power_up = "low";

dffeas \lpp_count_offset[4] (
	.clk(clk),
	.d(\Add1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~0_combout ),
	.q(\lpp_count_offset[4]~q ),
	.prn(vcc));
defparam \lpp_count_offset[4] .is_wysiwyg = "true";
defparam \lpp_count_offset[4] .power_up = "low";

dffeas fft_dirn_held_o(
	.clk(clk),
	.d(\fft_dirn_held_o~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_dirn_held_o~q ),
	.prn(vcc));
defparam fft_dirn_held_o.is_wysiwyg = "true";
defparam fft_dirn_held_o.power_up = "low";

dffeas \lpp_count[0] (
	.clk(clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_count[0]~q ),
	.prn(vcc));
defparam \lpp_count[0] .is_wysiwyg = "true";
defparam \lpp_count[0] .power_up = "low";

dffeas \lpp_count[1] (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_count[1]~q ),
	.prn(vcc));
defparam \lpp_count[1] .is_wysiwyg = "true";
defparam \lpp_count[1] .power_up = "low";

dffeas \lpp_count[2] (
	.clk(clk),
	.d(\lpp_count~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_count[2]~q ),
	.prn(vcc));
defparam \lpp_count[2] .is_wysiwyg = "true";
defparam \lpp_count[2] .power_up = "low";

dffeas \lpp_count[3] (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_count[3]~q ),
	.prn(vcc));
defparam \lpp_count[3] .is_wysiwyg = "true";
defparam \lpp_count[3] .power_up = "low";

dffeas \lpp_count[4] (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_count[4]~q ),
	.prn(vcc));
defparam \lpp_count[4] .is_wysiwyg = "true";
defparam \lpp_count[4] .power_up = "low";

dffeas \lpp_count[5] (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_count[5]~q ),
	.prn(vcc));
defparam \lpp_count[5] .is_wysiwyg = "true";
defparam \lpp_count[5] .power_up = "low";

dffeas fft_dirn_held(
	.clk(clk),
	.d(\fft_dirn~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_dirn_held~q ),
	.prn(vcc));
defparam fft_dirn_held.is_wysiwyg = "true";
defparam fft_dirn_held.power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lpp_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h00000000000000FF;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lpp_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h00000000000000FF;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lpp_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h00000000000000FF;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lpp_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h00000000000000FF;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lpp_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h00000000000000FF;
defparam \Add2~17 .shared_arith = "off";

cyclonev_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lpp_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h00000000000000FF;
defparam \Add2~21 .shared_arith = "off";

dffeas fft_dirn(
	.clk(clk),
	.d(\fft_dirn~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_dirn~q ),
	.prn(vcc));
defparam fft_dirn.is_wysiwyg = "true";
defparam fft_dirn.power_up = "low";

dffeas \data_rdy_vec[4] (
	.clk(clk),
	.d(\data_rdy_vec[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[4]~q ),
	.prn(vcc));
defparam \data_rdy_vec[4] .is_wysiwyg = "true";
defparam \data_rdy_vec[4] .power_up = "low";

dffeas \data_rdy_vec[3] (
	.clk(clk),
	.d(\data_rdy_vec[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[3]~q ),
	.prn(vcc));
defparam \data_rdy_vec[3] .is_wysiwyg = "true";
defparam \data_rdy_vec[3] .power_up = "low";

dffeas \data_rdy_vec[2] (
	.clk(clk),
	.d(\data_rdy_vec[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[2]~q ),
	.prn(vcc));
defparam \data_rdy_vec[2] .is_wysiwyg = "true";
defparam \data_rdy_vec[2] .power_up = "low";

dffeas \data_rdy_vec[1] (
	.clk(clk),
	.d(\data_rdy_vec[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[1]~q ),
	.prn(vcc));
defparam \data_rdy_vec[1] .is_wysiwyg = "true";
defparam \data_rdy_vec[1] .power_up = "low";

dffeas \data_rdy_vec[0] (
	.clk(clk),
	.d(\writer|data_rdy_int~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[0]~q ),
	.prn(vcc));
defparam \data_rdy_vec[0] .is_wysiwyg = "true";
defparam \data_rdy_vec[0] .power_up = "low";

dffeas \lpp_ram_data_out[3][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][10] .power_up = "low";

dffeas \lpp_ram_data_out[0][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][10] .power_up = "low";

dffeas \lpp_ram_data_out[1][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][10] .power_up = "low";

dffeas \lpp_ram_data_out[2][10] (
	.clk(clk),
	.d(\lpp_ram_data_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][10]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][10] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][10] .power_up = "low";

dffeas \lpp_ram_data_out[3][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][2] .power_up = "low";

dffeas \lpp_ram_data_out[0][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][2] .power_up = "low";

dffeas \lpp_ram_data_out[1][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][2] .power_up = "low";

dffeas \lpp_ram_data_out[2][2] (
	.clk(clk),
	.d(\lpp_ram_data_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][2]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][2] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][2] .power_up = "low";

dffeas \lpp_ram_data_out[3][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][11] .power_up = "low";

dffeas \lpp_ram_data_out[0][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][11] .power_up = "low";

dffeas \lpp_ram_data_out[1][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][11] .power_up = "low";

dffeas \lpp_ram_data_out[2][11] (
	.clk(clk),
	.d(\lpp_ram_data_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][11]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][11] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][11] .power_up = "low";

dffeas \lpp_ram_data_out[3][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][3] .power_up = "low";

dffeas \lpp_ram_data_out[0][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][3] .power_up = "low";

dffeas \lpp_ram_data_out[1][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][3] .power_up = "low";

dffeas \lpp_ram_data_out[2][3] (
	.clk(clk),
	.d(\lpp_ram_data_out~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][3]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][3] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][3] .power_up = "low";

dffeas \lpp_ram_data_out[3][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][12] .power_up = "low";

dffeas \lpp_ram_data_out[0][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][12] .power_up = "low";

dffeas \lpp_ram_data_out[1][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][12] .power_up = "low";

dffeas \lpp_ram_data_out[2][12] (
	.clk(clk),
	.d(\lpp_ram_data_out~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][12]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][12] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][12] .power_up = "low";

dffeas \lpp_ram_data_out[3][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][4] .power_up = "low";

dffeas \lpp_ram_data_out[0][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][4] .power_up = "low";

dffeas \lpp_ram_data_out[1][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][4] .power_up = "low";

dffeas \lpp_ram_data_out[2][4] (
	.clk(clk),
	.d(\lpp_ram_data_out~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][4]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][4] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][4] .power_up = "low";

dffeas \lpp_ram_data_out[3][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][13] .power_up = "low";

dffeas \lpp_ram_data_out[0][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][13] .power_up = "low";

dffeas \lpp_ram_data_out[1][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][13] .power_up = "low";

dffeas \lpp_ram_data_out[2][13] (
	.clk(clk),
	.d(\lpp_ram_data_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][13]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][13] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][13] .power_up = "low";

dffeas \lpp_ram_data_out[3][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][5] .power_up = "low";

dffeas \lpp_ram_data_out[0][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][5] .power_up = "low";

dffeas \lpp_ram_data_out[1][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][5] .power_up = "low";

dffeas \lpp_ram_data_out[2][5] (
	.clk(clk),
	.d(\lpp_ram_data_out~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][5]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][5] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][5] .power_up = "low";

dffeas \lpp_ram_data_out[3][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][14] .power_up = "low";

dffeas \lpp_ram_data_out[0][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][14] .power_up = "low";

dffeas \lpp_ram_data_out[1][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][14] .power_up = "low";

dffeas \lpp_ram_data_out[2][14] (
	.clk(clk),
	.d(\lpp_ram_data_out~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][14]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][14] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][14] .power_up = "low";

dffeas \lpp_ram_data_out[3][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][6] .power_up = "low";

dffeas \lpp_ram_data_out[0][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][6] .power_up = "low";

dffeas \lpp_ram_data_out[1][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][6] .power_up = "low";

dffeas \lpp_ram_data_out[2][6] (
	.clk(clk),
	.d(\lpp_ram_data_out~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][6]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][6] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][6] .power_up = "low";

dffeas \lpp_ram_data_out[3][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][15] .power_up = "low";

dffeas \lpp_ram_data_out[0][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][15] .power_up = "low";

dffeas \lpp_ram_data_out[1][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][15] .power_up = "low";

dffeas \lpp_ram_data_out[2][15] (
	.clk(clk),
	.d(\lpp_ram_data_out~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][15]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][15] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][15] .power_up = "low";

dffeas \lpp_ram_data_out[3][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][7] .power_up = "low";

dffeas \lpp_ram_data_out[0][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][7] .power_up = "low";

dffeas \lpp_ram_data_out[1][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][7] .power_up = "low";

dffeas \lpp_ram_data_out[2][7] (
	.clk(clk),
	.d(\lpp_ram_data_out~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][7]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][7] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][7] .power_up = "low";

dffeas lpp_sel(
	.clk(clk),
	.d(\lpp_sel~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_sel~q ),
	.prn(vcc));
defparam lpp_sel.is_wysiwyg = "true";
defparam lpp_sel.power_up = "low";

dffeas \lpp_ram_data_out[3][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][9] .power_up = "low";

dffeas \lpp_ram_data_out[0][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][9] .power_up = "low";

dffeas \lpp_ram_data_out[1][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][9] .power_up = "low";

dffeas \lpp_ram_data_out[2][9] (
	.clk(clk),
	.d(\lpp_ram_data_out~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][9]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][9] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][9] .power_up = "low";

dffeas \lpp_ram_data_out[3][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][1] .power_up = "low";

dffeas \lpp_ram_data_out[0][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][1] .power_up = "low";

dffeas \lpp_ram_data_out[1][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][1] .power_up = "low";

dffeas \lpp_ram_data_out[2][1] (
	.clk(clk),
	.d(\lpp_ram_data_out~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][1]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][1] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][1] .power_up = "low";

dffeas \wc_vec[3] (
	.clk(clk),
	.d(\wc_vec[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wc_vec[3]~q ),
	.prn(vcc));
defparam \wc_vec[3] .is_wysiwyg = "true";
defparam \wc_vec[3] .power_up = "low";

dffeas \rdaddress_c_bus[0] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[0]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[0] .power_up = "low";

dffeas \rdaddress_c_bus[13] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[13]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[13] .power_up = "low";

dffeas \rdaddress_c_bus[10] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[10]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[10] .power_up = "low";

dffeas \rdaddress_c_bus[3] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[3][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[3]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[3] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[3] .power_up = "low";

dffeas \wd_vec[3] (
	.clk(clk),
	.d(\wd_vec[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wd_vec[3]~q ),
	.prn(vcc));
defparam \wd_vec[3] .is_wysiwyg = "true";
defparam \wd_vec[3] .power_up = "low";

dffeas \rdaddress_c_bus[14] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[1][2]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[14]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[14] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[14] .power_up = "low";

dffeas \rdaddress_c_bus[15] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[15]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[15] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[15] .power_up = "low";

dffeas \rdaddress_c_bus[11] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[3][3]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[11]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[11] .power_up = "low";

dffeas \rdaddress_c_bus[7] (
	.clk(clk),
	.d(\gen_radix_4_last_pass:gen_M4K_output_sel:ram_cxb_rd_lpp|ram_in_reg[0][3]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\rdaddress_c_bus[7]~q ),
	.prn(vcc));
defparam \rdaddress_c_bus[7] .is_wysiwyg = "true";
defparam \rdaddress_c_bus[7] .power_up = "low";

dffeas \lpp_ram_data_out[3][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][8] .power_up = "low";

dffeas \lpp_ram_data_out[0][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][8] .power_up = "low";

dffeas \lpp_ram_data_out[1][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][8] .power_up = "low";

dffeas \lpp_ram_data_out[2][8] (
	.clk(clk),
	.d(\lpp_ram_data_out~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][8]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][8] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][8] .power_up = "low";

dffeas \lpp_ram_data_out[3][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[3][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[3][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[3][0] .power_up = "low";

dffeas \lpp_ram_data_out[0][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[0][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[0][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[0][0] .power_up = "low";

dffeas \lpp_ram_data_out[1][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[1][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[1][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[1][0] .power_up = "low";

dffeas \lpp_ram_data_out[2][0] (
	.clk(clk),
	.d(\lpp_ram_data_out~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\lpp_ram_data_out[2][0]~q ),
	.prn(vcc));
defparam \lpp_ram_data_out[2][0] .is_wysiwyg = "true";
defparam \lpp_ram_data_out[2][0] .power_up = "low";

dffeas \wc_vec[2] (
	.clk(clk),
	.d(\wc_vec[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wc_vec[2]~q ),
	.prn(vcc));
defparam \wc_vec[2] .is_wysiwyg = "true";
defparam \wc_vec[2] .power_up = "low";

dffeas \wd_vec[2] (
	.clk(clk),
	.d(\wd_vec[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wd_vec[2]~q ),
	.prn(vcc));
defparam \wd_vec[2] .is_wysiwyg = "true";
defparam \wd_vec[2] .power_up = "low";

dffeas \wc_vec[1] (
	.clk(clk),
	.d(\wc_vec[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wc_vec[1]~q ),
	.prn(vcc));
defparam \wc_vec[1] .is_wysiwyg = "true";
defparam \wc_vec[1] .power_up = "low";

dffeas \wd_vec[1] (
	.clk(clk),
	.d(\wd_vec[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wd_vec[1]~q ),
	.prn(vcc));
defparam \wd_vec[1] .is_wysiwyg = "true";
defparam \wd_vec[1] .power_up = "low";

dffeas \wc_vec[0] (
	.clk(clk),
	.d(\sel_we|wc_i~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wc_vec[0]~q ),
	.prn(vcc));
defparam \wc_vec[0] .is_wysiwyg = "true";
defparam \wc_vec[0] .power_up = "low";

dffeas \wd_vec[0] (
	.clk(clk),
	.d(\sel_we|wd_i~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wd_vec[0]~q ),
	.prn(vcc));
defparam \wd_vec[0] .is_wysiwyg = "true";
defparam \wd_vec[0] .power_up = "low";

dffeas \twiddle_data[0][1][0] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][0] .power_up = "low";

dffeas \twiddle_data[0][1][1] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][1] .power_up = "low";

dffeas \twiddle_data[0][1][2] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][2] .power_up = "low";

dffeas \twiddle_data[0][1][3] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][3] .power_up = "low";

dffeas \twiddle_data[0][1][4] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][4] .power_up = "low";

dffeas \twiddle_data[0][1][5] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][5] .power_up = "low";

dffeas \twiddle_data[0][1][6] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][6] .power_up = "low";

dffeas \twiddle_data[0][1][7] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[0][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[0][1][7] .power_up = "low";

dffeas \twiddle_data[0][0][7] (
	.clk(clk),
	.d(\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][7] .power_up = "low";

dffeas \twiddle_data[1][0][7] (
	.clk(clk),
	.d(\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][7] .power_up = "low";

dffeas \twiddle_data[1][1][0] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][0] .power_up = "low";

dffeas \twiddle_data[1][1][1] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][1] .power_up = "low";

dffeas \twiddle_data[1][1][2] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][2] .power_up = "low";

dffeas \twiddle_data[1][1][3] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][3] .power_up = "low";

dffeas \twiddle_data[1][1][4] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][4] .power_up = "low";

dffeas \twiddle_data[1][1][5] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][5] .power_up = "low";

dffeas \twiddle_data[1][1][6] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][6] .power_up = "low";

dffeas \twiddle_data[1][1][7] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[1][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[1][1][7] .power_up = "low";

dffeas \twiddle_data[2][0][7] (
	.clk(clk),
	.d(\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][7]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][7] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][7] .power_up = "low";

dffeas \twiddle_data[2][1][0] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][0]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][0] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][0] .power_up = "low";

dffeas \twiddle_data[2][1][1] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][1]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][1] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][1] .power_up = "low";

dffeas \twiddle_data[2][1][2] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][2]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][2] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][2] .power_up = "low";

dffeas \twiddle_data[2][1][3] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][3]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][3] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][3] .power_up = "low";

dffeas \twiddle_data[2][1][4] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][4]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][4] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][4] .power_up = "low";

dffeas \twiddle_data[2][1][5] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][5]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][5] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][5] .power_up = "low";

dffeas \twiddle_data[2][1][6] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][6]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][6] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][6] .power_up = "low";

dffeas \twiddle_data[2][1][7] (
	.clk(clk),
	.d(\twrom|gen_M4K:sin_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][1][7]~q ),
	.prn(vcc));
defparam \twiddle_data[2][1][7] .is_wysiwyg = "true";
defparam \twiddle_data[2][1][7] .power_up = "low";

dffeas \data_rdy_vec[10] (
	.clk(clk),
	.d(\data_rdy_vec[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[10]~q ),
	.prn(vcc));
defparam \data_rdy_vec[10] .is_wysiwyg = "true";
defparam \data_rdy_vec[10] .power_up = "low";

dffeas \data_rdy_vec[9] (
	.clk(clk),
	.d(\data_rdy_vec[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[9]~q ),
	.prn(vcc));
defparam \data_rdy_vec[9] .is_wysiwyg = "true";
defparam \data_rdy_vec[9] .power_up = "low";

dffeas \wren_b[1] (
	.clk(clk),
	.d(\wren_b~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_b[1]~q ),
	.prn(vcc));
defparam \wren_b[1] .is_wysiwyg = "true";
defparam \wren_b[1] .power_up = "low";

dffeas \wren_a[1] (
	.clk(clk),
	.d(\wren_a~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_a[1]~q ),
	.prn(vcc));
defparam \wren_a[1] .is_wysiwyg = "true";
defparam \wren_a[1] .power_up = "low";

dffeas \wren_b[2] (
	.clk(clk),
	.d(\wren_b~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_b[2]~q ),
	.prn(vcc));
defparam \wren_b[2] .is_wysiwyg = "true";
defparam \wren_b[2] .power_up = "low";

dffeas \wren_a[2] (
	.clk(clk),
	.d(\wren_a~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_a[2]~q ),
	.prn(vcc));
defparam \wren_a[2] .is_wysiwyg = "true";
defparam \wren_a[2] .power_up = "low";

dffeas \wren_b[3] (
	.clk(clk),
	.d(\wren_b~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_b[3]~q ),
	.prn(vcc));
defparam \wren_b[3] .is_wysiwyg = "true";
defparam \wren_b[3] .power_up = "low";

dffeas \wren_a[3] (
	.clk(clk),
	.d(\wren_a~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_a[3]~q ),
	.prn(vcc));
defparam \wren_a[3] .is_wysiwyg = "true";
defparam \wren_a[3] .power_up = "low";

dffeas \wren_b[0] (
	.clk(clk),
	.d(\wren_b~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_b[0]~q ),
	.prn(vcc));
defparam \wren_b[0] .is_wysiwyg = "true";
defparam \wren_b[0] .power_up = "low";

dffeas \wren_a[0] (
	.clk(clk),
	.d(\wren_a~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(!\global_clock_enable~0_combout ),
	.q(\wren_a[0]~q ),
	.prn(vcc));
defparam \wren_a[0] .is_wysiwyg = "true";
defparam \wren_a[0] .power_up = "low";

dffeas \data_rdy_vec[8] (
	.clk(clk),
	.d(\data_rdy_vec[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[8]~q ),
	.prn(vcc));
defparam \data_rdy_vec[8] .is_wysiwyg = "true";
defparam \data_rdy_vec[8] .power_up = "low";

dffeas \data_rdy_vec[7] (
	.clk(clk),
	.d(\data_rdy_vec[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[7]~q ),
	.prn(vcc));
defparam \data_rdy_vec[7] .is_wysiwyg = "true";
defparam \data_rdy_vec[7] .power_up = "low";

dffeas \core_real_in[6] (
	.clk(clk),
	.d(\data_real_in_reg[6]~q ),
	.asdata(\data_imag_in_reg[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[6]~q ),
	.prn(vcc));
defparam \core_real_in[6] .is_wysiwyg = "true";
defparam \core_real_in[6] .power_up = "low";

dffeas \core_real_in[5] (
	.clk(clk),
	.d(\data_real_in_reg[5]~q ),
	.asdata(\data_imag_in_reg[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[5]~q ),
	.prn(vcc));
defparam \core_real_in[5] .is_wysiwyg = "true";
defparam \core_real_in[5] .power_up = "low";

dffeas \core_real_in[2] (
	.clk(clk),
	.d(\data_real_in_reg[2]~q ),
	.asdata(\data_imag_in_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[2]~q ),
	.prn(vcc));
defparam \core_real_in[2] .is_wysiwyg = "true";
defparam \core_real_in[2] .power_up = "low";

dffeas \core_real_in[3] (
	.clk(clk),
	.d(\data_real_in_reg[3]~q ),
	.asdata(\data_imag_in_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[3]~q ),
	.prn(vcc));
defparam \core_real_in[3] .is_wysiwyg = "true";
defparam \core_real_in[3] .power_up = "low";

dffeas \core_real_in[4] (
	.clk(clk),
	.d(\data_real_in_reg[4]~q ),
	.asdata(\data_imag_in_reg[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[4]~q ),
	.prn(vcc));
defparam \core_real_in[4] .is_wysiwyg = "true";
defparam \core_real_in[4] .power_up = "low";

dffeas \core_real_in[7] (
	.clk(clk),
	.d(\data_real_in_reg[7]~q ),
	.asdata(\data_imag_in_reg[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[7]~q ),
	.prn(vcc));
defparam \core_real_in[7] .is_wysiwyg = "true";
defparam \core_real_in[7] .power_up = "low";

dffeas \core_imag_in[7] (
	.clk(clk),
	.d(\data_imag_in_reg[7]~q ),
	.asdata(\data_real_in_reg[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[7]~q ),
	.prn(vcc));
defparam \core_imag_in[7] .is_wysiwyg = "true";
defparam \core_imag_in[7] .power_up = "low";

dffeas \core_imag_in[6] (
	.clk(clk),
	.d(\data_imag_in_reg[6]~q ),
	.asdata(\data_real_in_reg[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[6]~q ),
	.prn(vcc));
defparam \core_imag_in[6] .is_wysiwyg = "true";
defparam \core_imag_in[6] .power_up = "low";

dffeas \core_imag_in[3] (
	.clk(clk),
	.d(\data_imag_in_reg[3]~q ),
	.asdata(\data_real_in_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[3]~q ),
	.prn(vcc));
defparam \core_imag_in[3] .is_wysiwyg = "true";
defparam \core_imag_in[3] .power_up = "low";

dffeas \core_imag_in[4] (
	.clk(clk),
	.d(\data_imag_in_reg[4]~q ),
	.asdata(\data_real_in_reg[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[4]~q ),
	.prn(vcc));
defparam \core_imag_in[4] .is_wysiwyg = "true";
defparam \core_imag_in[4] .power_up = "low";

dffeas \core_imag_in[5] (
	.clk(clk),
	.d(\data_imag_in_reg[5]~q ),
	.asdata(\data_real_in_reg[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[5]~q ),
	.prn(vcc));
defparam \core_imag_in[5] .is_wysiwyg = "true";
defparam \core_imag_in[5] .power_up = "low";

dffeas \core_imag_in[2] (
	.clk(clk),
	.d(\data_imag_in_reg[2]~q ),
	.asdata(\data_real_in_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[2]~q ),
	.prn(vcc));
defparam \core_imag_in[2] .is_wysiwyg = "true";
defparam \core_imag_in[2] .power_up = "low";

dffeas \core_real_in[0] (
	.clk(clk),
	.d(\data_real_in_reg[0]~q ),
	.asdata(\data_imag_in_reg[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[0]~q ),
	.prn(vcc));
defparam \core_real_in[0] .is_wysiwyg = "true";
defparam \core_real_in[0] .power_up = "low";

dffeas \core_real_in[1] (
	.clk(clk),
	.d(\data_real_in_reg[1]~q ),
	.asdata(\data_imag_in_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_real_in[1]~q ),
	.prn(vcc));
defparam \core_real_in[1] .is_wysiwyg = "true";
defparam \core_real_in[1] .power_up = "low";

dffeas \core_imag_in[0] (
	.clk(clk),
	.d(\data_imag_in_reg[0]~q ),
	.asdata(\data_real_in_reg[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[0]~q ),
	.prn(vcc));
defparam \core_imag_in[0] .is_wysiwyg = "true";
defparam \core_imag_in[0] .power_up = "low";

dffeas \core_imag_in[1] (
	.clk(clk),
	.d(\data_imag_in_reg[1]~q ),
	.asdata(\data_real_in_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(\fft_dirn~q ),
	.ena(!\global_clock_enable~0_combout ),
	.q(\core_imag_in[1]~q ),
	.prn(vcc));
defparam \core_imag_in[1] .is_wysiwyg = "true";
defparam \core_imag_in[1] .power_up = "low";

dffeas \data_rdy_vec[6] (
	.clk(clk),
	.d(\data_rdy_vec[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[6]~q ),
	.prn(vcc));
defparam \data_rdy_vec[6] .is_wysiwyg = "true";
defparam \data_rdy_vec[6] .power_up = "low";

dffeas \data_real_in_reg[6] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[6]~q ),
	.prn(vcc));
defparam \data_real_in_reg[6] .is_wysiwyg = "true";
defparam \data_real_in_reg[6] .power_up = "low";

dffeas \data_imag_in_reg[6] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[6]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[6] .is_wysiwyg = "true";
defparam \data_imag_in_reg[6] .power_up = "low";

dffeas \data_real_in_reg[5] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[5]~q ),
	.prn(vcc));
defparam \data_real_in_reg[5] .is_wysiwyg = "true";
defparam \data_real_in_reg[5] .power_up = "low";

dffeas \data_imag_in_reg[5] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[5]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[5] .is_wysiwyg = "true";
defparam \data_imag_in_reg[5] .power_up = "low";

dffeas \data_real_in_reg[2] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[2]~q ),
	.prn(vcc));
defparam \data_real_in_reg[2] .is_wysiwyg = "true";
defparam \data_real_in_reg[2] .power_up = "low";

dffeas \data_imag_in_reg[2] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[2]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[2] .is_wysiwyg = "true";
defparam \data_imag_in_reg[2] .power_up = "low";

dffeas \data_real_in_reg[3] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[3]~q ),
	.prn(vcc));
defparam \data_real_in_reg[3] .is_wysiwyg = "true";
defparam \data_real_in_reg[3] .power_up = "low";

dffeas \data_imag_in_reg[3] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[3]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[3] .is_wysiwyg = "true";
defparam \data_imag_in_reg[3] .power_up = "low";

dffeas \data_real_in_reg[4] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[4]~q ),
	.prn(vcc));
defparam \data_real_in_reg[4] .is_wysiwyg = "true";
defparam \data_real_in_reg[4] .power_up = "low";

dffeas \data_imag_in_reg[4] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[4]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[4] .is_wysiwyg = "true";
defparam \data_imag_in_reg[4] .power_up = "low";

dffeas \data_real_in_reg[7] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[7]~q ),
	.prn(vcc));
defparam \data_real_in_reg[7] .is_wysiwyg = "true";
defparam \data_real_in_reg[7] .power_up = "low";

dffeas \data_imag_in_reg[7] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[7]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[7] .is_wysiwyg = "true";
defparam \data_imag_in_reg[7] .power_up = "low";

dffeas \data_real_in_reg[0] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[0]~q ),
	.prn(vcc));
defparam \data_real_in_reg[0] .is_wysiwyg = "true";
defparam \data_real_in_reg[0] .power_up = "low";

dffeas \data_imag_in_reg[0] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[0]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[0] .is_wysiwyg = "true";
defparam \data_imag_in_reg[0] .power_up = "low";

dffeas \data_real_in_reg[1] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_real_in_reg[1]~q ),
	.prn(vcc));
defparam \data_real_in_reg[1] .is_wysiwyg = "true";
defparam \data_real_in_reg[1] .power_up = "low";

dffeas \data_imag_in_reg[1] (
	.clk(clk),
	.d(\auk_dsp_atlantic_sink_1|normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_imag_in_reg[1]~q ),
	.prn(vcc));
defparam \data_imag_in_reg[1] .is_wysiwyg = "true";
defparam \data_imag_in_reg[1] .power_up = "low";

dffeas \data_rdy_vec[5] (
	.clk(clk),
	.d(\data_rdy_vec[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_rdy_vec[5]~q ),
	.prn(vcc));
defparam \data_rdy_vec[5] .is_wysiwyg = "true";
defparam \data_rdy_vec[5] .power_up = "low";

cyclonev_lcell_comb \data_count_sig[2]~5 (
	.dataa(!\data_count_sig[0]~q ),
	.datab(!\master_source_sop~q ),
	.datac(!\LessThan0~1_combout ),
	.datad(!\global_clock_enable~0_combout ),
	.datae(!\data_sample_counter~0_combout ),
	.dataf(!\data_count_sig[2]~q ),
	.datag(!\data_count_sig[1]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_count_sig[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_count_sig[2]~5 .extended_lut = "on";
defparam \data_count_sig[2]~5 .lut_mask = 64'hB77BF7FBB77BF7FB;
defparam \data_count_sig[2]~5 .shared_arith = "off";

dffeas master_sink_ena(
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\master_sink_ena~q ),
	.prn(vcc));
defparam master_sink_ena.is_wysiwyg = "true";
defparam master_sink_ena.power_up = "low";

dffeas sink_ready_ctrl_d(
	.clk(clk),
	.d(\auk_dsp_interface_controller_1|sink_ready_ctrl~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_ready_ctrl_d~q ),
	.prn(vcc));
defparam sink_ready_ctrl_d.is_wysiwyg = "true";
defparam sink_ready_ctrl_d.power_up = "low";

dffeas sop(
	.clk(clk),
	.d(\sop~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sop~q ),
	.prn(vcc));
defparam sop.is_wysiwyg = "true";
defparam sop.power_up = "low";

dffeas \data_count_sig[3] (
	.clk(clk),
	.d(\data_count_sig[3]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_count_sig[3]~q ),
	.prn(vcc));
defparam \data_count_sig[3] .is_wysiwyg = "true";
defparam \data_count_sig[3] .power_up = "low";

dffeas \data_count_sig[2] (
	.clk(clk),
	.d(\data_count_sig[2]~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_count_sig[2]~q ),
	.prn(vcc));
defparam \data_count_sig[2] .is_wysiwyg = "true";
defparam \data_count_sig[2] .power_up = "low";

dffeas \data_count_sig[1] (
	.clk(clk),
	.d(\data_count_sig[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_count_sig[1]~q ),
	.prn(vcc));
defparam \data_count_sig[1] .is_wysiwyg = "true";
defparam \data_count_sig[1] .power_up = "low";

dffeas \data_count_sig[0] (
	.clk(clk),
	.d(\data_count_sig~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\data_count_sig[0]~q ),
	.prn(vcc));
defparam \data_count_sig[0] .is_wysiwyg = "true";
defparam \data_count_sig[0] .power_up = "low";

dffeas \data_count_sig[5] (
	.clk(clk),
	.d(\data_count_sig[5]~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_count_sig[5]~q ),
	.prn(vcc));
defparam \data_count_sig[5] .is_wysiwyg = "true";
defparam \data_count_sig[5] .power_up = "low";

dffeas \data_count_sig[4] (
	.clk(clk),
	.d(\data_count_sig[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\data_count_sig[4]~q ),
	.prn(vcc));
defparam \data_count_sig[4] .is_wysiwyg = "true";
defparam \data_count_sig[4] .power_up = "low";

dffeas \exponent_out[0] (
	.clk(clk),
	.d(\exponent_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\exponent_out[0]~q ),
	.prn(vcc));
defparam \exponent_out[0] .is_wysiwyg = "true";
defparam \exponent_out[0] .power_up = "low";

dffeas \exponent_out[1] (
	.clk(clk),
	.d(\exponent_out~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\exponent_out[1]~q ),
	.prn(vcc));
defparam \exponent_out[1] .is_wysiwyg = "true";
defparam \exponent_out[1] .power_up = "low";

dffeas \exponent_out[2] (
	.clk(clk),
	.d(\exponent_out~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\exponent_out[2]~q ),
	.prn(vcc));
defparam \exponent_out[2] .is_wysiwyg = "true";
defparam \exponent_out[2] .power_up = "low";

dffeas \exponent_out[3] (
	.clk(clk),
	.d(\exponent_out~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\exponent_out[3]~q ),
	.prn(vcc));
defparam \exponent_out[3] .is_wysiwyg = "true";
defparam \exponent_out[3] .power_up = "low";

dffeas \exponent_out[4] (
	.clk(clk),
	.d(\exponent_out~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\exponent_out[4]~q ),
	.prn(vcc));
defparam \exponent_out[4] .is_wysiwyg = "true";
defparam \exponent_out[4] .power_up = "low";

dffeas \exponent_out[5] (
	.clk(clk),
	.d(\exponent_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\exponent_out[5]~q ),
	.prn(vcc));
defparam \exponent_out[5] .is_wysiwyg = "true";
defparam \exponent_out[5] .power_up = "low";

cyclonev_lcell_comb \global_clock_enable~0 (
	.dataa(!\sink_ready_ctrl_d~q ),
	.datab(!\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datac(!\sop~q ),
	.datad(!\auk_dsp_atlantic_source_1|source_stall_int_d~q ),
	.datae(!\auk_dsp_interface_controller_1|stall_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\global_clock_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \global_clock_enable~0 .extended_lut = "off";
defparam \global_clock_enable~0 .lut_mask = 64'hFFFF96FFFFFF96FF;
defparam \global_clock_enable~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_in_work~0 (
	.dataa(!\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.datab(!\sink_in_work~q ),
	.datac(!\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_in_work~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_in_work~0 .extended_lut = "off";
defparam \sink_in_work~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \sink_in_work~0 .shared_arith = "off";

cyclonev_lcell_comb \sop~0 (
	.dataa(!\auk_dsp_atlantic_sink_1|send_eop_s~q ),
	.datab(!\sink_ready_ctrl_d~q ),
	.datac(!\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datad(!\sop~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop~0 .extended_lut = "off";
defparam \sop~0 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \sop~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\data_count_sig[2]~q ),
	.datab(!\data_count_sig[1]~q ),
	.datac(!\data_count_sig[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\data_count_sig[4]~q ),
	.datab(!\data_count_sig[3]~q ),
	.datac(!\data_count_sig[2]~q ),
	.datad(!\data_count_sig[1]~q ),
	.datae(!\data_count_sig[0]~q ),
	.dataf(!\data_count_sig[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \data_sample_counter~0 (
	.dataa(!\data_count_sig[4]~q ),
	.datab(!\data_count_sig[3]~q ),
	.datac(!\data_count_sig[2]~q ),
	.datad(!\data_count_sig[1]~q ),
	.datae(!\data_count_sig[0]~q ),
	.dataf(!\data_count_sig[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_sample_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_sample_counter~0 .extended_lut = "off";
defparam \data_sample_counter~0 .lut_mask = 64'h6996966996696996;
defparam \data_sample_counter~0 .shared_arith = "off";

dffeas master_source_sop(
	.clk(clk),
	.d(\master_source_sop~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\master_source_sop~q ),
	.prn(vcc));
defparam master_source_sop.is_wysiwyg = "true";
defparam master_source_sop.power_up = "low";

cyclonev_lcell_comb \data_count_sig[3]~0 (
	.dataa(!\data_count_sig[3]~q ),
	.datab(!\global_clock_enable~0_combout ),
	.datac(!\LessThan0~0_combout ),
	.datad(!\LessThan0~1_combout ),
	.datae(!\data_sample_counter~0_combout ),
	.dataf(!\master_source_sop~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_count_sig[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_count_sig[3]~0 .extended_lut = "off";
defparam \data_count_sig[3]~0 .lut_mask = 64'hFFFFFFFF69FF96FF;
defparam \data_count_sig[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \data_count_sig[1]~1 (
	.dataa(!\data_count_sig[1]~q ),
	.datab(!\data_count_sig[0]~q ),
	.datac(!\global_clock_enable~0_combout ),
	.datad(!\LessThan0~1_combout ),
	.datae(!\data_sample_counter~0_combout ),
	.dataf(!\master_source_sop~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_count_sig[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_count_sig[1]~1 .extended_lut = "off";
defparam \data_count_sig[1]~1 .lut_mask = 64'hFFFFFFFF69FF96FF;
defparam \data_count_sig[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \data_count_sig~2 (
	.dataa(!\data_count_sig[0]~q ),
	.datab(!\data_sample_counter~0_combout ),
	.datac(!\master_source_sop~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_count_sig~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_count_sig~2 .extended_lut = "off";
defparam \data_count_sig~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \data_count_sig~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!\data_count_sig[3]~q ),
	.datab(!\data_count_sig[2]~q ),
	.datac(!\data_count_sig[1]~q ),
	.datad(!\data_count_sig[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~2 .shared_arith = "off";

cyclonev_lcell_comb \data_count_sig[5]~3 (
	.dataa(!\data_count_sig[4]~q ),
	.datab(!\data_count_sig[5]~q ),
	.datac(!\global_clock_enable~0_combout ),
	.datad(!\LessThan0~2_combout ),
	.datae(!\data_sample_counter~0_combout ),
	.dataf(!\master_source_sop~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_count_sig[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_count_sig[5]~3 .extended_lut = "off";
defparam \data_count_sig[5]~3 .lut_mask = 64'hFFFFFFFFFFFF6996;
defparam \data_count_sig[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \data_count_sig[4]~4 (
	.dataa(!\data_count_sig[4]~q ),
	.datab(!\data_count_sig[5]~q ),
	.datac(!\global_clock_enable~0_combout ),
	.datad(!\LessThan0~2_combout ),
	.datae(!\data_sample_counter~0_combout ),
	.dataf(!\master_source_sop~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_count_sig[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_count_sig[4]~4 .extended_lut = "off";
defparam \data_count_sig[4]~4 .lut_mask = 64'hFFFFFFFFDEEDEDDE;
defparam \data_count_sig[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \fft_imag_out[1]~0 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_imag_out[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_imag_out[1]~0 .extended_lut = "off";
defparam \fft_imag_out[1]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \fft_imag_out[1]~0 .shared_arith = "off";

dffeas \blk_exp_accum[0] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[0]~q ),
	.prn(vcc));
defparam \blk_exp_accum[0] .is_wysiwyg = "true";
defparam \blk_exp_accum[0] .power_up = "low";

cyclonev_lcell_comb \exponent_out~0 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\blk_exp_accum[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\exponent_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \exponent_out~0 .extended_lut = "off";
defparam \exponent_out~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \exponent_out~0 .shared_arith = "off";

dffeas \blk_exp_accum[1] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[1]~q ),
	.prn(vcc));
defparam \blk_exp_accum[1] .is_wysiwyg = "true";
defparam \blk_exp_accum[1] .power_up = "low";

cyclonev_lcell_comb \exponent_out~1 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\blk_exp_accum[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\exponent_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \exponent_out~1 .extended_lut = "off";
defparam \exponent_out~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \exponent_out~1 .shared_arith = "off";

dffeas \blk_exp_accum[2] (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[2]~q ),
	.prn(vcc));
defparam \blk_exp_accum[2] .is_wysiwyg = "true";
defparam \blk_exp_accum[2] .power_up = "low";

cyclonev_lcell_comb \exponent_out~2 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\blk_exp_accum[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\exponent_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \exponent_out~2 .extended_lut = "off";
defparam \exponent_out~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \exponent_out~2 .shared_arith = "off";

dffeas \blk_exp_accum[3] (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[3]~q ),
	.prn(vcc));
defparam \blk_exp_accum[3] .is_wysiwyg = "true";
defparam \blk_exp_accum[3] .power_up = "low";

cyclonev_lcell_comb \exponent_out~3 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\blk_exp_accum[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\exponent_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \exponent_out~3 .extended_lut = "off";
defparam \exponent_out~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \exponent_out~3 .shared_arith = "off";

dffeas \blk_exp_accum[4] (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[4]~q ),
	.prn(vcc));
defparam \blk_exp_accum[4] .is_wysiwyg = "true";
defparam \blk_exp_accum[4] .power_up = "low";

cyclonev_lcell_comb \exponent_out~4 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\blk_exp_accum[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\exponent_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \exponent_out~4 .extended_lut = "off";
defparam \exponent_out~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \exponent_out~4 .shared_arith = "off";

dffeas \blk_exp_accum[5] (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\blk_exp_accum[5]~q ),
	.prn(vcc));
defparam \blk_exp_accum[5] .is_wysiwyg = "true";
defparam \blk_exp_accum[5] .power_up = "low";

cyclonev_lcell_comb \exponent_out~5 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\blk_exp_accum[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\exponent_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \exponent_out~5 .extended_lut = "off";
defparam \exponent_out~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \exponent_out~5 .shared_arith = "off";

dffeas \fft_s2_cur.IDLE (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s2_cur.IDLE~1_combout ),
	.q(\fft_s2_cur.IDLE~q ),
	.prn(vcc));
defparam \fft_s2_cur.IDLE .is_wysiwyg = "true";
defparam \fft_s2_cur.IDLE .power_up = "low";

cyclonev_lcell_comb WideNor1(
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam WideNor1.shared_arith = "off";

cyclonev_lcell_comb \master_source_sop~0 (
	.dataa(!reset_n),
	.datab(!\oe~q ),
	.datac(!\sop_out~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_source_sop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_source_sop~0 .extended_lut = "off";
defparam \master_source_sop~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \master_source_sop~0 .shared_arith = "off";

dffeas \fft_s2_cur.FIRST_LPP_C (
	.clk(clk),
	.d(\fft_s2_cur~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\fft_s2_cur.FIRST_LPP_C~q ),
	.prn(vcc));
defparam \fft_s2_cur.FIRST_LPP_C .is_wysiwyg = "true";
defparam \fft_s2_cur.FIRST_LPP_C .power_up = "low";

cyclonev_lcell_comb \fft_dirn_stream~0 (
	.dataa(!\fft_dirn_stream~q ),
	.datab(!\fft_dirn_held_o2~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_dirn_stream~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_dirn_stream~0 .extended_lut = "off";
defparam \fft_dirn_stream~0 .lut_mask = 64'h5353535353535353;
defparam \fft_dirn_stream~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!\blk_exp_accum[0]~q ),
	.datab(!\fft_s2_cur.IDLE~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\gen_dft_1:bfpc|blk_exp[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!\blk_exp_accum[1]~q ),
	.datab(!\fft_s2_cur.IDLE~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\gen_dft_1:bfpc|blk_exp[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\blk_exp_accum[2]~q ),
	.datab(!\fft_s2_cur.IDLE~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\gen_dft_1:bfpc|blk_exp[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\blk_exp_accum[3]~q ),
	.datab(!\fft_s2_cur.IDLE~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\gen_dft_1:bfpc|blk_exp[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\blk_exp_accum[4]~q ),
	.datab(!\fft_s2_cur.IDLE~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\gen_dft_1:bfpc|blk_exp[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\blk_exp_accum[5]~q ),
	.datab(!\fft_s2_cur.IDLE~q ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\gen_dft_1:bfpc|blk_exp[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \Selector0~0 .shared_arith = "off";

dffeas \fft_s2_cur.LPP_C_OUTPUT (
	.clk(clk),
	.d(\fft_s2_cur.LPP_C_OUTPUT~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fft_s2_cur.LPP_C_OUTPUT~q ),
	.prn(vcc));
defparam \fft_s2_cur.LPP_C_OUTPUT .is_wysiwyg = "true";
defparam \fft_s2_cur.LPP_C_OUTPUT .power_up = "low";

dffeas \lpp_count_offset[0] (
	.clk(clk),
	.d(\lpp_count_offset~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\lpp_count_offset[0]~0_combout ),
	.q(\lpp_count_offset[0]~q ),
	.prn(vcc));
defparam \lpp_count_offset[0] .is_wysiwyg = "true";
defparam \lpp_count_offset[0] .power_up = "low";

cyclonev_lcell_comb \fft_s2_cur.IDLE~0 (
	.dataa(!\lpp_count_offset[0]~q ),
	.datab(!\lpp_count_offset[1]~q ),
	.datac(!\lpp_count_offset[2]~q ),
	.datad(!\lpp_count_offset[3]~q ),
	.datae(!\lpp_count_offset[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_s2_cur.IDLE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_s2_cur.IDLE~0 .extended_lut = "off";
defparam \fft_s2_cur.IDLE~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \fft_s2_cur.IDLE~0 .shared_arith = "off";

cyclonev_lcell_comb \fft_s2_cur.IDLE~1 (
	.dataa(!reset_n),
	.datab(!\global_clock_enable~0_combout ),
	.datac(!\fft_s2_cur.LPP_C_OUTPUT~q ),
	.datad(!\lpp_count_offset[5]~q ),
	.datae(!\fft_s2_cur.IDLE~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_s2_cur.IDLE~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_s2_cur.IDLE~1 .extended_lut = "off";
defparam \fft_s2_cur.IDLE~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \fft_s2_cur.IDLE~1 .shared_arith = "off";

dffeas \fft_s2_cur.LAST_LPP_C (
	.clk(clk),
	.d(\fft_s2_cur.LAST_LPP_C~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fft_s2_cur.IDLE~1_combout ),
	.q(\fft_s2_cur.LAST_LPP_C~q ),
	.prn(vcc));
defparam \fft_s2_cur.LAST_LPP_C .is_wysiwyg = "true";
defparam \fft_s2_cur.LAST_LPP_C .power_up = "low";

cyclonev_lcell_comb \Selector17~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\delay_lpp_en|tdl_arr[5]~q ),
	.datad(!\fft_s2_cur.LAST_LPP_C~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector17~0 .extended_lut = "off";
defparam \Selector17~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \Selector17~0 .shared_arith = "off";

cyclonev_lcell_comb \fft_dirn_held_o2~0 (
	.dataa(!\fft_dirn_held_o2~q ),
	.datab(!\fft_dirn_held_o~q ),
	.datac(!\gen_le256_mk:ctrl|blk_done_int~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_dirn_held_o2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_dirn_held_o2~0 .extended_lut = "off";
defparam \fft_dirn_held_o2~0 .lut_mask = 64'h5353535353535353;
defparam \fft_dirn_held_o2~0 .shared_arith = "off";

cyclonev_lcell_comb \fft_s2_cur~9 (
	.dataa(!reset_n),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\delay_lpp_en|tdl_arr[5]~q ),
	.datad(!\fft_s2_cur.LAST_LPP_C~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_s2_cur~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_s2_cur~9 .extended_lut = "off";
defparam \fft_s2_cur~9 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \fft_s2_cur~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_s2_cur.LPP_C_OUTPUT~0 (
	.dataa(!reset_n),
	.datab(!\global_clock_enable~0_combout ),
	.datac(!\fft_s2_cur.FIRST_LPP_C~q ),
	.datad(!\fft_s2_cur.LPP_C_OUTPUT~q ),
	.datae(!\lpp_count_offset[5]~q ),
	.dataf(!\fft_s2_cur.IDLE~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_s2_cur.LPP_C_OUTPUT~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_s2_cur.LPP_C_OUTPUT~0 .extended_lut = "off";
defparam \fft_s2_cur.LPP_C_OUTPUT~0 .lut_mask = 64'hFFFF7FFFDFFF5FFF;
defparam \fft_s2_cur.LPP_C_OUTPUT~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\lpp_count[0]~q ),
	.datab(!\lpp_count[1]~q ),
	.datac(!\lpp_count[2]~q ),
	.datad(!\lpp_count[3]~q ),
	.datae(!\lpp_count[4]~q ),
	.dataf(!\lpp_count[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h6996966996696996;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \lpp_count_offset[0]~0 (
	.dataa(!reset_n),
	.datab(!\global_clock_enable~0_combout ),
	.datac(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_count_offset[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_count_offset[0]~0 .extended_lut = "off";
defparam \lpp_count_offset[0]~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \lpp_count_offset[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \lpp_count_offset~1 (
	.dataa(!reset_n),
	.datab(!\lpp_count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_count_offset~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_count_offset~1 .extended_lut = "off";
defparam \lpp_count_offset~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \lpp_count_offset~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\lpp_count[0]~q ),
	.datab(!\lpp_count[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6666666666666666;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~2 (
	.dataa(!\lpp_count[0]~q ),
	.datab(!\lpp_count[1]~q ),
	.datac(!\lpp_count[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~2 .extended_lut = "off";
defparam \Add1~2 .lut_mask = 64'h9696969696969696;
defparam \Add1~2 .shared_arith = "off";

cyclonev_lcell_comb \Add1~3 (
	.dataa(!\lpp_count[0]~q ),
	.datab(!\lpp_count[1]~q ),
	.datac(!\lpp_count[2]~q ),
	.datad(!\lpp_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~3 .extended_lut = "off";
defparam \Add1~3 .lut_mask = 64'h6996699669966996;
defparam \Add1~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~4 (
	.dataa(!\lpp_count[0]~q ),
	.datab(!\lpp_count[1]~q ),
	.datac(!\lpp_count[2]~q ),
	.datad(!\lpp_count[3]~q ),
	.datae(!\lpp_count[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~4 .extended_lut = "off";
defparam \Add1~4 .lut_mask = 64'h9669699696696996;
defparam \Add1~4 .shared_arith = "off";

cyclonev_lcell_comb \fft_s2_cur.LAST_LPP_C~0 (
	.dataa(!reset_n),
	.datab(!\fft_s2_cur.LPP_C_OUTPUT~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_s2_cur.LAST_LPP_C~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_s2_cur.LAST_LPP_C~0 .extended_lut = "off";
defparam \fft_s2_cur.LAST_LPP_C~0 .lut_mask = 64'h7777777777777777;
defparam \fft_s2_cur.LAST_LPP_C~0 .shared_arith = "off";

cyclonev_lcell_comb \fft_dirn_held_o~0 (
	.dataa(!\fft_dirn_held_o~q ),
	.datab(!\writer|next_block~q ),
	.datac(!\fft_dirn_held~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_dirn_held_o~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_dirn_held_o~0 .extended_lut = "off";
defparam \fft_dirn_held_o~0 .lut_mask = 64'h4747474747474747;
defparam \fft_dirn_held_o~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector11~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\Add2~1_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector11~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\Add2~5_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector10~0 .shared_arith = "off";

cyclonev_lcell_comb \lpp_count~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\Add2~9_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_count~0 .extended_lut = "off";
defparam \lpp_count~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \lpp_count~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\Add2~13_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector9~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\Add2~17_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!\fft_s2_cur.IDLE~q ),
	.datab(!\fft_s2_cur.WAIT_FOR_LPP_INPUT~q ),
	.datac(!\Add2~21_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector7~0 .shared_arith = "off";

dffeas inv_i(
	.clk(clk),
	.d(\inv_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\inv_i~q ),
	.prn(vcc));
defparam inv_i.is_wysiwyg = "true";
defparam inv_i.power_up = "low";

cyclonev_lcell_comb \fft_dirn~0 (
	.dataa(!\auk_dsp_atlantic_sink_1|send_sop_s~q ),
	.datab(!\fft_dirn~q ),
	.datac(!\inv_i~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fft_dirn~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fft_dirn~0 .extended_lut = "off";
defparam \fft_dirn~0 .lut_mask = 64'h2727272727272727;
defparam \fft_dirn~0 .shared_arith = "off";

cyclonev_lcell_comb \inv_i~0 (
	.dataa(!sink_valid),
	.datab(!\inv_i~q ),
	.datac(!inverse_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\inv_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \inv_i~0 .extended_lut = "off";
defparam \inv_i~0 .lut_mask = 64'h2727272727272727;
defparam \inv_i~0 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~0 (
	.dataa(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datab(!\lpp_sel~q ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~0 .extended_lut = "off";
defparam \lpp_ram_data_out~0 .lut_mask = 64'h4747474747474747;
defparam \lpp_ram_data_out~0 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~1 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~1 .extended_lut = "off";
defparam \lpp_ram_data_out~1 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~1 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~2 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~2 .extended_lut = "off";
defparam \lpp_ram_data_out~2 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~2 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~3 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~3 .extended_lut = "off";
defparam \lpp_ram_data_out~3 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~3 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~4 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~4 .extended_lut = "off";
defparam \lpp_ram_data_out~4 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~4 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~5 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~5 .extended_lut = "off";
defparam \lpp_ram_data_out~5 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~5 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~6 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~6 .extended_lut = "off";
defparam \lpp_ram_data_out~6 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~6 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~7 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~7 .extended_lut = "off";
defparam \lpp_ram_data_out~7 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~7 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~8 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~8 .extended_lut = "off";
defparam \lpp_ram_data_out~8 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~8 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~9 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~9 .extended_lut = "off";
defparam \lpp_ram_data_out~9 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~9 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~10 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~10 .extended_lut = "off";
defparam \lpp_ram_data_out~10 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~10 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~11 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~11 .extended_lut = "off";
defparam \lpp_ram_data_out~11 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~11 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~12 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~12 .extended_lut = "off";
defparam \lpp_ram_data_out~12 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~12 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~13 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~13 .extended_lut = "off";
defparam \lpp_ram_data_out~13 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~13 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~14 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~14 .extended_lut = "off";
defparam \lpp_ram_data_out~14 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~14 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~15 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~15 .extended_lut = "off";
defparam \lpp_ram_data_out~15 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~15 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~16 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~16 .extended_lut = "off";
defparam \lpp_ram_data_out~16 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~16 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~17 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~17 .extended_lut = "off";
defparam \lpp_ram_data_out~17 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~17 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~18 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~18 .extended_lut = "off";
defparam \lpp_ram_data_out~18 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~18 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~19 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~19 .extended_lut = "off";
defparam \lpp_ram_data_out~19 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~19 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~20 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~20 .extended_lut = "off";
defparam \lpp_ram_data_out~20 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~20 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~21 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~21 .extended_lut = "off";
defparam \lpp_ram_data_out~21 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~21 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~22 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~22 .extended_lut = "off";
defparam \lpp_ram_data_out~22 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~22 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~23 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~23 .extended_lut = "off";
defparam \lpp_ram_data_out~23 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~23 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~24 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~24 .extended_lut = "off";
defparam \lpp_ram_data_out~24 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~24 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~25 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~25 .extended_lut = "off";
defparam \lpp_ram_data_out~25 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~25 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~26 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~26 .extended_lut = "off";
defparam \lpp_ram_data_out~26 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~26 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~27 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~27 .extended_lut = "off";
defparam \lpp_ram_data_out~27 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~27 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~28 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~28 .extended_lut = "off";
defparam \lpp_ram_data_out~28 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~28 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~29 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~29 .extended_lut = "off";
defparam \lpp_ram_data_out~29 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~29 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~30 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~30 .extended_lut = "off";
defparam \lpp_ram_data_out~30 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~30 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~31 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~31 .extended_lut = "off";
defparam \lpp_ram_data_out~31 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~31 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~32 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~32 .extended_lut = "off";
defparam \lpp_ram_data_out~32 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~32 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~33 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~33 .extended_lut = "off";
defparam \lpp_ram_data_out~33 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~33 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~34 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~34 .extended_lut = "off";
defparam \lpp_ram_data_out~34 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~34 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~35 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~35 .extended_lut = "off";
defparam \lpp_ram_data_out~35 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~35 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~36 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~36 .extended_lut = "off";
defparam \lpp_ram_data_out~36 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~36 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~37 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~37 .extended_lut = "off";
defparam \lpp_ram_data_out~37 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~37 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~38 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~38 .extended_lut = "off";
defparam \lpp_ram_data_out~38 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~38 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~39 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~39 .extended_lut = "off";
defparam \lpp_ram_data_out~39 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~39 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~40 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~40 .extended_lut = "off";
defparam \lpp_ram_data_out~40 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~40 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~41 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~41 .extended_lut = "off";
defparam \lpp_ram_data_out~41 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~41 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~42 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~42 .extended_lut = "off";
defparam \lpp_ram_data_out~42 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~42 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~43 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~43 .extended_lut = "off";
defparam \lpp_ram_data_out~43 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~43 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~44 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~44 .extended_lut = "off";
defparam \lpp_ram_data_out~44 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~44 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~45 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~45 .extended_lut = "off";
defparam \lpp_ram_data_out~45 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~45 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~46 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~46 .extended_lut = "off";
defparam \lpp_ram_data_out~46 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~46 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~47 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~47 .extended_lut = "off";
defparam \lpp_ram_data_out~47 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~47 .shared_arith = "off";

cyclonev_lcell_comb \lpp_sel~0 (
	.dataa(!\gen_radix_4_last_pass:gen_lpp_addr|delay_en|tdl_arr[4]~q ),
	.datab(!\lpp_sel~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_sel~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_sel~0 .extended_lut = "off";
defparam \lpp_sel~0 .lut_mask = 64'h6666666666666666;
defparam \lpp_sel~0 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~48 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~48 .extended_lut = "off";
defparam \lpp_ram_data_out~48 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~48 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~49 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~49 .extended_lut = "off";
defparam \lpp_ram_data_out~49 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~49 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~50 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~50 .extended_lut = "off";
defparam \lpp_ram_data_out~50 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~50 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~51 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~51 .extended_lut = "off";
defparam \lpp_ram_data_out~51 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~51 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~52 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~52 .extended_lut = "off";
defparam \lpp_ram_data_out~52 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~52 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~53 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~53 .extended_lut = "off";
defparam \lpp_ram_data_out~53 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~53 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~54 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~54 .extended_lut = "off";
defparam \lpp_ram_data_out~54 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~54 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~55 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~55 .extended_lut = "off";
defparam \lpp_ram_data_out~55 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~55 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~56 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~56 .extended_lut = "off";
defparam \lpp_ram_data_out~56 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~56 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~57 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~57 .extended_lut = "off";
defparam \lpp_ram_data_out~57 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~57 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~58 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~58 .extended_lut = "off";
defparam \lpp_ram_data_out~58 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~58 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~59 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~59 .extended_lut = "off";
defparam \lpp_ram_data_out~59 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~59 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~60 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:3:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~60 .extended_lut = "off";
defparam \lpp_ram_data_out~60 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~60 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~61 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:0:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~61 .extended_lut = "off";
defparam \lpp_ram_data_out~61 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~61 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~62 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:1:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~62 .extended_lut = "off";
defparam \lpp_ram_data_out~62 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~62 .shared_arith = "off";

cyclonev_lcell_comb \lpp_ram_data_out~63 (
	.dataa(!\lpp_sel~q ),
	.datab(!\gen_M4K_Output:dat_C|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datac(!\gen_M4K_Output:dat_D|gen_rams:2:dat_A|gen_M4K:ram_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lpp_ram_data_out~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lpp_ram_data_out~63 .extended_lut = "off";
defparam \lpp_ram_data_out~63 .lut_mask = 64'h2727272727272727;
defparam \lpp_ram_data_out~63 .shared_arith = "off";

dffeas en_slb(
	.clk(clk),
	.d(\en_slb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\en_slb~q ),
	.prn(vcc));
defparam en_slb.is_wysiwyg = "true";
defparam en_slb.power_up = "low";

dffeas \p_tdl[0][0] (
	.clk(clk),
	.d(\gen_le256_mk:ctrl|p[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[0][0]~q ),
	.prn(vcc));
defparam \p_tdl[0][0] .is_wysiwyg = "true";
defparam \p_tdl[0][0] .power_up = "low";

dffeas \p_tdl[0][1] (
	.clk(clk),
	.d(\gen_le256_mk:ctrl|p[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[0][1]~q ),
	.prn(vcc));
defparam \p_tdl[0][1] .is_wysiwyg = "true";
defparam \p_tdl[0][1] .power_up = "low";

cyclonev_lcell_comb \en_slb~0 (
	.dataa(!\gen_le256_mk:ctrl|p[1]~q ),
	.datab(!\gen_le256_mk:ctrl|p[0]~q ),
	.datac(!\delay_ctrl_np|tdl_arr[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\en_slb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \en_slb~0 .extended_lut = "off";
defparam \en_slb~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \en_slb~0 .shared_arith = "off";

dffeas \ram_a_not_b_vec[26] (
	.clk(clk),
	.d(\ram_a_not_b_vec~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[26]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[26] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[26] .power_up = "low";

dffeas \p_cd_en[0] (
	.clk(clk),
	.d(\p_tdl[12][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_cd_en[0]~q ),
	.prn(vcc));
defparam \p_cd_en[0] .is_wysiwyg = "true";
defparam \p_cd_en[0] .power_up = "low";

dffeas \p_cd_en[1] (
	.clk(clk),
	.d(\p_tdl[12][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_cd_en[1]~q ),
	.prn(vcc));
defparam \p_cd_en[1] .is_wysiwyg = "true";
defparam \p_cd_en[1] .power_up = "low";

dffeas \twiddle_data[0][0][0] (
	.clk(clk),
	.d(\twiddle_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][0] .power_up = "low";

dffeas \twiddle_data[0][0][1] (
	.clk(clk),
	.d(\twiddle_data~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][1] .power_up = "low";

dffeas \twiddle_data[0][0][2] (
	.clk(clk),
	.d(\twiddle_data~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][2] .power_up = "low";

dffeas \twiddle_data[0][0][3] (
	.clk(clk),
	.d(\twiddle_data~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][3] .power_up = "low";

dffeas \twiddle_data[0][0][4] (
	.clk(clk),
	.d(\twiddle_data~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][4] .power_up = "low";

dffeas \twiddle_data[0][0][5] (
	.clk(clk),
	.d(\twiddle_data~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][5] .power_up = "low";

dffeas \twiddle_data[0][0][6] (
	.clk(clk),
	.d(\twiddle_data~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[0][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[0][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[0][0][6] .power_up = "low";

dffeas \twiddle_data[1][0][0] (
	.clk(clk),
	.d(\twiddle_data~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][0] .power_up = "low";

dffeas \twiddle_data[1][0][1] (
	.clk(clk),
	.d(\twiddle_data~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][1] .power_up = "low";

dffeas \twiddle_data[1][0][2] (
	.clk(clk),
	.d(\twiddle_data~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][2] .power_up = "low";

dffeas \twiddle_data[1][0][3] (
	.clk(clk),
	.d(\twiddle_data~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][3] .power_up = "low";

dffeas \twiddle_data[1][0][4] (
	.clk(clk),
	.d(\twiddle_data~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][4] .power_up = "low";

dffeas \twiddle_data[1][0][5] (
	.clk(clk),
	.d(\twiddle_data~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][5] .power_up = "low";

dffeas \twiddle_data[1][0][6] (
	.clk(clk),
	.d(\twiddle_data~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[1][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[1][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[1][0][6] .power_up = "low";

dffeas \twiddle_data[2][0][0] (
	.clk(clk),
	.d(\twiddle_data~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][0]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][0] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][0] .power_up = "low";

dffeas \twiddle_data[2][0][1] (
	.clk(clk),
	.d(\twiddle_data~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][1]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][1] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][1] .power_up = "low";

dffeas \twiddle_data[2][0][2] (
	.clk(clk),
	.d(\twiddle_data~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][2]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][2] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][2] .power_up = "low";

dffeas \twiddle_data[2][0][3] (
	.clk(clk),
	.d(\twiddle_data~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][3]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][3] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][3] .power_up = "low";

dffeas \twiddle_data[2][0][4] (
	.clk(clk),
	.d(\twiddle_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][4]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][4] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][4] .power_up = "low";

dffeas \twiddle_data[2][0][5] (
	.clk(clk),
	.d(\twiddle_data~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][5]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][5] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][5] .power_up = "low";

dffeas \twiddle_data[2][0][6] (
	.clk(clk),
	.d(\twiddle_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\twiddle_data[2][0][6]~q ),
	.prn(vcc));
defparam \twiddle_data[2][0][6] .is_wysiwyg = "true";
defparam \twiddle_data[2][0][6] .power_up = "low";

dffeas \ram_a_not_b_vec[25] (
	.clk(clk),
	.d(\ram_a_not_b_vec~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[25]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[25] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[25] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~0 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~0 .extended_lut = "off";
defparam \ram_a_not_b_vec~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~0 .shared_arith = "off";

dffeas \p_tdl[12][0] (
	.clk(clk),
	.d(\p_tdl[11][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[12][0]~q ),
	.prn(vcc));
defparam \p_tdl[12][0] .is_wysiwyg = "true";
defparam \p_tdl[12][0] .power_up = "low";

dffeas \p_tdl[12][1] (
	.clk(clk),
	.d(\p_tdl[11][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[12][1]~q ),
	.prn(vcc));
defparam \p_tdl[12][1] .is_wysiwyg = "true";
defparam \p_tdl[12][1] .power_up = "low";

cyclonev_lcell_comb \twiddle_data~0 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~0 .extended_lut = "off";
defparam \twiddle_data~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~0 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~1 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~1 .extended_lut = "off";
defparam \twiddle_data~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~1 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~2 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~2 .extended_lut = "off";
defparam \twiddle_data~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~2 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~3 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~3 .extended_lut = "off";
defparam \twiddle_data~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~3 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~4 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~4 .extended_lut = "off";
defparam \twiddle_data~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~4 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~5 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~5 .extended_lut = "off";
defparam \twiddle_data~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~5 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~6 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_1n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~6 .extended_lut = "off";
defparam \twiddle_data~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~6 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~7 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~7 .extended_lut = "off";
defparam \twiddle_data~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~7 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~8 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~8 .extended_lut = "off";
defparam \twiddle_data~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~8 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~9 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~9 .extended_lut = "off";
defparam \twiddle_data~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~9 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~10 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~10 .extended_lut = "off";
defparam \twiddle_data~10 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~10 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~11 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~11 .extended_lut = "off";
defparam \twiddle_data~11 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~11 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~12 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~12 .extended_lut = "off";
defparam \twiddle_data~12 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~12 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~13 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_2n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~13 .extended_lut = "off";
defparam \twiddle_data~13 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~13 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~14 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~14 .extended_lut = "off";
defparam \twiddle_data~14 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~14 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~15 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~15 .extended_lut = "off";
defparam \twiddle_data~15 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~15 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~16 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~16 .extended_lut = "off";
defparam \twiddle_data~16 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~16 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~17 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~17 .extended_lut = "off";
defparam \twiddle_data~17 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~17 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~18 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~18 .extended_lut = "off";
defparam \twiddle_data~18 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~18 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~19 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~19 .extended_lut = "off";
defparam \twiddle_data~19 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~19 .shared_arith = "off";

cyclonev_lcell_comb \twiddle_data~20 (
	.dataa(!reset_n),
	.datab(!\twrom|gen_M4K:cos_3n|gen_auto:rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\twiddle_data~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \twiddle_data~20 .extended_lut = "off";
defparam \twiddle_data~20 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \twiddle_data~20 .shared_arith = "off";

dffeas \ram_a_not_b_vec[24] (
	.clk(clk),
	.d(\ram_a_not_b_vec~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[24]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[24] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[24] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~1 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~1 .extended_lut = "off";
defparam \ram_a_not_b_vec~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~1 .shared_arith = "off";

dffeas \p_tdl[11][0] (
	.clk(clk),
	.d(\p_tdl[10][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[11][0]~q ),
	.prn(vcc));
defparam \p_tdl[11][0] .is_wysiwyg = "true";
defparam \p_tdl[11][0] .power_up = "low";

dffeas \p_tdl[11][1] (
	.clk(clk),
	.d(\p_tdl[10][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[11][1]~q ),
	.prn(vcc));
defparam \p_tdl[11][1] .is_wysiwyg = "true";
defparam \p_tdl[11][1] .power_up = "low";

dffeas \ram_a_not_b_vec[23] (
	.clk(clk),
	.d(\ram_a_not_b_vec~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[23]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[23] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[23] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~2 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~2 .extended_lut = "off";
defparam \ram_a_not_b_vec~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~2 .shared_arith = "off";

dffeas \p_tdl[10][0] (
	.clk(clk),
	.d(\p_tdl[9][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[10][0]~q ),
	.prn(vcc));
defparam \p_tdl[10][0] .is_wysiwyg = "true";
defparam \p_tdl[10][0] .power_up = "low";

dffeas \p_tdl[10][1] (
	.clk(clk),
	.d(\p_tdl[9][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[10][1]~q ),
	.prn(vcc));
defparam \p_tdl[10][1] .is_wysiwyg = "true";
defparam \p_tdl[10][1] .power_up = "low";

dffeas \ram_a_not_b_vec[22] (
	.clk(clk),
	.d(\ram_a_not_b_vec~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[22]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[22] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[22] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~3 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~3 .extended_lut = "off";
defparam \ram_a_not_b_vec~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~3 .shared_arith = "off";

dffeas \p_tdl[9][0] (
	.clk(clk),
	.d(\p_tdl[8][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[9][0]~q ),
	.prn(vcc));
defparam \p_tdl[9][0] .is_wysiwyg = "true";
defparam \p_tdl[9][0] .power_up = "low";

dffeas \p_tdl[9][1] (
	.clk(clk),
	.d(\p_tdl[8][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[9][1]~q ),
	.prn(vcc));
defparam \p_tdl[9][1] .is_wysiwyg = "true";
defparam \p_tdl[9][1] .power_up = "low";

dffeas \ram_a_not_b_vec[21] (
	.clk(clk),
	.d(\ram_a_not_b_vec~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[21]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[21] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[21] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~4 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~4 .extended_lut = "off";
defparam \ram_a_not_b_vec~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~4 .shared_arith = "off";

dffeas \p_tdl[8][0] (
	.clk(clk),
	.d(\p_tdl[7][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[8][0]~q ),
	.prn(vcc));
defparam \p_tdl[8][0] .is_wysiwyg = "true";
defparam \p_tdl[8][0] .power_up = "low";

dffeas \p_tdl[8][1] (
	.clk(clk),
	.d(\p_tdl[7][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[8][1]~q ),
	.prn(vcc));
defparam \p_tdl[8][1] .is_wysiwyg = "true";
defparam \p_tdl[8][1] .power_up = "low";

dffeas \ram_a_not_b_vec[20] (
	.clk(clk),
	.d(\ram_a_not_b_vec~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[20]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[20] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[20] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~5 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~5 .extended_lut = "off";
defparam \ram_a_not_b_vec~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~5 .shared_arith = "off";

dffeas \p_tdl[7][0] (
	.clk(clk),
	.d(\p_tdl[6][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[7][0]~q ),
	.prn(vcc));
defparam \p_tdl[7][0] .is_wysiwyg = "true";
defparam \p_tdl[7][0] .power_up = "low";

dffeas \p_tdl[7][1] (
	.clk(clk),
	.d(\p_tdl[6][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[7][1]~q ),
	.prn(vcc));
defparam \p_tdl[7][1] .is_wysiwyg = "true";
defparam \p_tdl[7][1] .power_up = "low";

dffeas \ram_a_not_b_vec[19] (
	.clk(clk),
	.d(\ram_a_not_b_vec~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[19]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[19] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[19] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~6 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~6 .extended_lut = "off";
defparam \ram_a_not_b_vec~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~6 .shared_arith = "off";

dffeas \p_tdl[6][0] (
	.clk(clk),
	.d(\p_tdl[5][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[6][0]~q ),
	.prn(vcc));
defparam \p_tdl[6][0] .is_wysiwyg = "true";
defparam \p_tdl[6][0] .power_up = "low";

dffeas \p_tdl[6][1] (
	.clk(clk),
	.d(\p_tdl[5][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[6][1]~q ),
	.prn(vcc));
defparam \p_tdl[6][1] .is_wysiwyg = "true";
defparam \p_tdl[6][1] .power_up = "low";

dffeas \sw_r_tdl[4][0] (
	.clk(clk),
	.d(\sw_r_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[4][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[4][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[4][0] .power_up = "low";

dffeas \sw_r_tdl[4][1] (
	.clk(clk),
	.d(\sw_r_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[4][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[4][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[4][1] .power_up = "low";

dffeas \ram_a_not_b_vec[18] (
	.clk(clk),
	.d(\ram_a_not_b_vec~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[18]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[18] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[18] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~7 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~7 .extended_lut = "off";
defparam \ram_a_not_b_vec~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~7 .shared_arith = "off";

dffeas \p_tdl[5][0] (
	.clk(clk),
	.d(\p_tdl[4][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[5][0]~q ),
	.prn(vcc));
defparam \p_tdl[5][0] .is_wysiwyg = "true";
defparam \p_tdl[5][0] .power_up = "low";

dffeas \p_tdl[5][1] (
	.clk(clk),
	.d(\p_tdl[4][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[5][1]~q ),
	.prn(vcc));
defparam \p_tdl[5][1] .is_wysiwyg = "true";
defparam \p_tdl[5][1] .power_up = "low";

dffeas \ram_a_not_b_vec[10] (
	.clk(clk),
	.d(\ram_a_not_b_vec~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[10]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[10] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[10] .power_up = "low";

dffeas \sw_r_tdl[3][0] (
	.clk(clk),
	.d(\sw_r_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[3][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[3][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[3][0] .power_up = "low";

dffeas \sw_r_tdl[3][1] (
	.clk(clk),
	.d(\sw_r_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[3][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[3][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[3][1] .power_up = "low";

dffeas \ram_a_not_b_vec[17] (
	.clk(clk),
	.d(\ram_a_not_b_vec~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[17]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[17] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[17] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~8 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~8 .extended_lut = "off";
defparam \ram_a_not_b_vec~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~8 .shared_arith = "off";

dffeas \p_tdl[4][0] (
	.clk(clk),
	.d(\p_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[4][0]~q ),
	.prn(vcc));
defparam \p_tdl[4][0] .is_wysiwyg = "true";
defparam \p_tdl[4][0] .power_up = "low";

dffeas \p_tdl[4][1] (
	.clk(clk),
	.d(\p_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[4][1]~q ),
	.prn(vcc));
defparam \p_tdl[4][1] .is_wysiwyg = "true";
defparam \p_tdl[4][1] .power_up = "low";

dffeas \ram_a_not_b_vec[9] (
	.clk(clk),
	.d(\ram_a_not_b_vec~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[9]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[9] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[9] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~9 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~9 .extended_lut = "off";
defparam \ram_a_not_b_vec~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~9 .shared_arith = "off";

dffeas \sw_r_tdl[2][0] (
	.clk(clk),
	.d(\sw_r_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[2][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[2][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[2][0] .power_up = "low";

dffeas \sw_r_tdl[2][1] (
	.clk(clk),
	.d(\sw_r_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[2][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[2][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[2][1] .power_up = "low";

dffeas \ram_a_not_b_vec[16] (
	.clk(clk),
	.d(\ram_a_not_b_vec~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[16]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[16] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[16] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~10 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~10 .extended_lut = "off";
defparam \ram_a_not_b_vec~10 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~10 .shared_arith = "off";

dffeas \p_tdl[3][0] (
	.clk(clk),
	.d(\p_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[3][0]~q ),
	.prn(vcc));
defparam \p_tdl[3][0] .is_wysiwyg = "true";
defparam \p_tdl[3][0] .power_up = "low";

dffeas \p_tdl[3][1] (
	.clk(clk),
	.d(\p_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[3][1]~q ),
	.prn(vcc));
defparam \p_tdl[3][1] .is_wysiwyg = "true";
defparam \p_tdl[3][1] .power_up = "low";

dffeas \ram_a_not_b_vec[8] (
	.clk(clk),
	.d(\ram_a_not_b_vec~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[8]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[8] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[8] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~11 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~11 .extended_lut = "off";
defparam \ram_a_not_b_vec~11 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~11 .shared_arith = "off";

dffeas \ram_a_not_b_vec[1] (
	.clk(clk),
	.d(\ram_a_not_b_vec~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[1]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[1] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[1] .power_up = "low";

cyclonev_lcell_comb \wren_b~0 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_b~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_b~0 .extended_lut = "off";
defparam \wren_b~0 .lut_mask = 64'h4747474747474747;
defparam \wren_b~0 .shared_arith = "off";

dffeas \ram_a_not_b_vec[7] (
	.clk(clk),
	.d(\ram_a_not_b_vec~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[7]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[7] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[7] .power_up = "low";

cyclonev_lcell_comb sel_anb_addr(
	.dataa(!\data_rdy_vec[10]~q ),
	.datab(!\ram_a_not_b_vec[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sel_anb_addr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam sel_anb_addr.extended_lut = "off";
defparam sel_anb_addr.lut_mask = 64'h7777777777777777;
defparam sel_anb_addr.shared_arith = "off";

cyclonev_lcell_comb \wren_a~0 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_a~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_a~0 .extended_lut = "off";
defparam \wren_a~0 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \wren_a~0 .shared_arith = "off";

cyclonev_lcell_comb \wren_b~1 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_b~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_b~1 .extended_lut = "off";
defparam \wren_b~1 .lut_mask = 64'h4747474747474747;
defparam \wren_b~1 .shared_arith = "off";

cyclonev_lcell_comb \wren_a~1 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_a~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_a~1 .extended_lut = "off";
defparam \wren_a~1 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \wren_a~1 .shared_arith = "off";

cyclonev_lcell_comb \wren_b~2 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_b~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_b~2 .extended_lut = "off";
defparam \wren_b~2 .lut_mask = 64'h4747474747474747;
defparam \wren_b~2 .shared_arith = "off";

cyclonev_lcell_comb \wren_a~2 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_a~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_a~2 .extended_lut = "off";
defparam \wren_a~2 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \wren_a~2 .shared_arith = "off";

cyclonev_lcell_comb \wren_b~3 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_b~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_b~3 .extended_lut = "off";
defparam \wren_b~3 .lut_mask = 64'h4747474747474747;
defparam \wren_b~3 .shared_arith = "off";

cyclonev_lcell_comb \wren_a~3 (
	.dataa(!\ram_a_not_b_vec[24]~q ),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(!\writer|wren[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren_a~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren_a~3 .extended_lut = "off";
defparam \wren_a~3 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \wren_a~3 .shared_arith = "off";

dffeas \sw_r_tdl[1][0] (
	.clk(clk),
	.d(\sw_r_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[1][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[1][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[1][0] .power_up = "low";

dffeas \sw_r_tdl[1][1] (
	.clk(clk),
	.d(\sw_r_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[1][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[1][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[1][1] .power_up = "low";

dffeas \ram_a_not_b_vec[15] (
	.clk(clk),
	.d(\ram_a_not_b_vec~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[15]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[15] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[15] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~12 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~12 .extended_lut = "off";
defparam \ram_a_not_b_vec~12 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~12 .shared_arith = "off";

dffeas \p_tdl[2][0] (
	.clk(clk),
	.d(\p_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[2][0]~q ),
	.prn(vcc));
defparam \p_tdl[2][0] .is_wysiwyg = "true";
defparam \p_tdl[2][0] .power_up = "low";

dffeas \p_tdl[2][1] (
	.clk(clk),
	.d(\p_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[2][1]~q ),
	.prn(vcc));
defparam \p_tdl[2][1] .is_wysiwyg = "true";
defparam \p_tdl[2][1] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~13 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~13 .extended_lut = "off";
defparam \ram_a_not_b_vec~13 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~13 .shared_arith = "off";

dffeas \ram_a_not_b_vec[0] (
	.clk(clk),
	.d(\ram_a_not_b_vec~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[0]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[0] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[0] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~14 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~14 .extended_lut = "off";
defparam \ram_a_not_b_vec~14 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~14 .shared_arith = "off";

dffeas \ram_a_not_b_vec[6] (
	.clk(clk),
	.d(\ram_a_not_b_vec~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[6]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[6] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[6] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~15 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~15 .extended_lut = "off";
defparam \ram_a_not_b_vec~15 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~15 .shared_arith = "off";

dffeas \sw_r_tdl[0][0] (
	.clk(clk),
	.d(\rd_adgen|sw[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[0][0]~q ),
	.prn(vcc));
defparam \sw_r_tdl[0][0] .is_wysiwyg = "true";
defparam \sw_r_tdl[0][0] .power_up = "low";

dffeas \sw_r_tdl[0][1] (
	.clk(clk),
	.d(\rd_adgen|sw[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\sw_r_tdl[0][1]~q ),
	.prn(vcc));
defparam \sw_r_tdl[0][1] .is_wysiwyg = "true";
defparam \sw_r_tdl[0][1] .power_up = "low";

dffeas \ram_a_not_b_vec[14] (
	.clk(clk),
	.d(\ram_a_not_b_vec~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[14]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[14] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[14] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~16 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~16 .extended_lut = "off";
defparam \ram_a_not_b_vec~16 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~16 .shared_arith = "off";

dffeas \p_tdl[1][0] (
	.clk(clk),
	.d(\p_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[1][0]~q ),
	.prn(vcc));
defparam \p_tdl[1][0] .is_wysiwyg = "true";
defparam \p_tdl[1][0] .power_up = "low";

dffeas \p_tdl[1][1] (
	.clk(clk),
	.d(\p_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\p_tdl[1][1]~q ),
	.prn(vcc));
defparam \p_tdl[1][1] .is_wysiwyg = "true";
defparam \p_tdl[1][1] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~17 (
	.dataa(!reset_n),
	.datab(!\writer|anb~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~17 .extended_lut = "off";
defparam \ram_a_not_b_vec~17 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~17 .shared_arith = "off";

dffeas \ram_a_not_b_vec[5] (
	.clk(clk),
	.d(\ram_a_not_b_vec~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[5]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[5] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[5] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~18 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~18 .extended_lut = "off";
defparam \ram_a_not_b_vec~18 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~18 .shared_arith = "off";

dffeas \ram_a_not_b_vec[13] (
	.clk(clk),
	.d(\ram_a_not_b_vec~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[13]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[13] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[13] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~19 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~19 .extended_lut = "off";
defparam \ram_a_not_b_vec~19 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~19 .shared_arith = "off";

dffeas \ram_a_not_b_vec[4] (
	.clk(clk),
	.d(\ram_a_not_b_vec~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[4]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[4] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[4] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~20 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~20 .extended_lut = "off";
defparam \ram_a_not_b_vec~20 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~20 .shared_arith = "off";

dffeas \ram_a_not_b_vec[12] (
	.clk(clk),
	.d(\ram_a_not_b_vec~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[12]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[12] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[12] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~21 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~21 .extended_lut = "off";
defparam \ram_a_not_b_vec~21 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~21 .shared_arith = "off";

dffeas \ram_a_not_b_vec[3] (
	.clk(clk),
	.d(\ram_a_not_b_vec~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[3]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[3] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[3] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~22 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~22 .extended_lut = "off";
defparam \ram_a_not_b_vec~22 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~22 .shared_arith = "off";

dffeas \ram_a_not_b_vec[11] (
	.clk(clk),
	.d(\ram_a_not_b_vec~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[11]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[11] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[11] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~23 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~23 .extended_lut = "off";
defparam \ram_a_not_b_vec~23 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~23 .shared_arith = "off";

dffeas \ram_a_not_b_vec[2] (
	.clk(clk),
	.d(\ram_a_not_b_vec~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\global_clock_enable~0_combout ),
	.q(\ram_a_not_b_vec[2]~q ),
	.prn(vcc));
defparam \ram_a_not_b_vec[2] .is_wysiwyg = "true";
defparam \ram_a_not_b_vec[2] .power_up = "low";

cyclonev_lcell_comb \ram_a_not_b_vec~24 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~24 .extended_lut = "off";
defparam \ram_a_not_b_vec~24 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~24 .shared_arith = "off";

cyclonev_lcell_comb \ram_a_not_b_vec~25 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~25 .extended_lut = "off";
defparam \ram_a_not_b_vec~25 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~25 .shared_arith = "off";

cyclonev_lcell_comb \ram_a_not_b_vec~26 (
	.dataa(!reset_n),
	.datab(!\ram_a_not_b_vec[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_a_not_b_vec~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_a_not_b_vec~26 .extended_lut = "off";
defparam \ram_a_not_b_vec~26 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ram_a_not_b_vec~26 .shared_arith = "off";

endmodule

module IFFT_asj_fft_3dp_rom (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	q_a_01,
	q_a_11,
	q_a_21,
	q_a_31,
	q_a_41,
	q_a_51,
	q_a_61,
	q_a_71,
	q_a_02,
	q_a_12,
	q_a_22,
	q_a_32,
	q_a_42,
	q_a_52,
	q_a_62,
	q_a_72,
	q_a_03,
	q_a_13,
	q_a_23,
	q_a_33,
	q_a_43,
	q_a_53,
	q_a_63,
	q_a_73,
	q_a_04,
	q_a_14,
	q_a_24,
	q_a_34,
	q_a_44,
	q_a_54,
	q_a_64,
	q_a_74,
	q_a_05,
	q_a_15,
	q_a_25,
	q_a_35,
	q_a_45,
	q_a_55,
	q_a_65,
	q_a_75,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
output 	q_a_01;
output 	q_a_11;
output 	q_a_21;
output 	q_a_31;
output 	q_a_41;
output 	q_a_51;
output 	q_a_61;
output 	q_a_71;
output 	q_a_02;
output 	q_a_12;
output 	q_a_22;
output 	q_a_32;
output 	q_a_42;
output 	q_a_52;
output 	q_a_62;
output 	q_a_72;
output 	q_a_03;
output 	q_a_13;
output 	q_a_23;
output 	q_a_33;
output 	q_a_43;
output 	q_a_53;
output 	q_a_63;
output 	q_a_73;
output 	q_a_04;
output 	q_a_14;
output 	q_a_24;
output 	q_a_34;
output 	q_a_44;
output 	q_a_54;
output 	q_a_64;
output 	q_a_74;
output 	q_a_05;
output 	q_a_15;
output 	q_a_25;
output 	q_a_35;
output 	q_a_45;
output 	q_a_55;
output 	q_a_65;
output 	q_a_75;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_twid_rom_2 \gen_M4K:cos_3n (
	.q_a_0(q_a_04),
	.q_a_1(q_a_14),
	.q_a_2(q_a_24),
	.q_a_3(q_a_34),
	.q_a_4(q_a_44),
	.q_a_5(q_a_54),
	.q_a_6(q_a_64),
	.q_a_7(q_a_74),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

IFFT_twid_rom_1 \gen_M4K:cos_2n (
	.q_a_0(q_a_02),
	.q_a_1(q_a_12),
	.q_a_2(q_a_22),
	.q_a_3(q_a_32),
	.q_a_4(q_a_42),
	.q_a_5(q_a_52),
	.q_a_6(q_a_62),
	.q_a_7(q_a_72),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

IFFT_twid_rom \gen_M4K:cos_1n (
	.q_a_0(q_a_01),
	.q_a_1(q_a_11),
	.q_a_2(q_a_21),
	.q_a_3(q_a_31),
	.q_a_4(q_a_41),
	.q_a_5(q_a_51),
	.q_a_6(q_a_61),
	.q_a_7(q_a_71),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

IFFT_twid_rom_5 \gen_M4K:sin_3n (
	.q_a_0(q_a_05),
	.q_a_1(q_a_15),
	.q_a_2(q_a_25),
	.q_a_3(q_a_35),
	.q_a_4(q_a_45),
	.q_a_5(q_a_55),
	.q_a_6(q_a_65),
	.q_a_7(q_a_75),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

IFFT_twid_rom_4 \gen_M4K:sin_2n (
	.q_a_0(q_a_03),
	.q_a_1(q_a_13),
	.q_a_2(q_a_23),
	.q_a_3(q_a_33),
	.q_a_4(q_a_43),
	.q_a_5(q_a_53),
	.q_a_6(q_a_63),
	.q_a_7(q_a_73),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

IFFT_twid_rom_3 \gen_M4K:sin_1n (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_twid_rom (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_single_port_rom \gen_auto:rom_component (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_single_port_rom (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_1 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_1 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_4e34 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_4e34 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "7615";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "05CB";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "AC17";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "C94F";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "5B3F";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "38FF";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "07FF";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "IFFT_fft_ii_0_1n64cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_4e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "0000";

endmodule

module IFFT_twid_rom_1 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_single_port_rom_1 \gen_auto:rom_component (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_single_port_rom_1 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_2 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_2 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_5e34 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_5e34 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "CEE7";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "F639";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "3627";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "4C9B";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "28D7";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "1A4F";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "063F";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "IFFT_fft_ii_0_2n64cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_5e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FE00";

endmodule

module IFFT_twid_rom_2 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_single_port_rom_2 \gen_auto:rom_component (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_single_port_rom_2 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_3 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_3 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_6e34 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_6e34 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "D459";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "BD47";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "21E1";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "F027";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "E21B";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "4157";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "80CF";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "IFFT_fft_ii_0_3n64cos.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:cos_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_6e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFC0";

endmodule

module IFFT_twid_rom_3 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_single_port_rom_3 \gen_auto:rom_component (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_single_port_rom_3 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_4 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_4 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_9e34 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_9e34 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "50DC";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "A740";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "D06A";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "E526";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "F9B4";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FE38";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFC0";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "IFFT_fft_ii_0_1n64sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_1n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_9e34:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "0000";

endmodule

module IFFT_twid_rom_4 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_single_port_rom_4 \gen_auto:rom_component (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_single_port_rom_4 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_5 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_5 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_ae34 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_ae34 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "E7CE";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "3938";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "27C8";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "9BB2";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "D7D6";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "4FE4";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "3FF8";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "IFFT_fft_ii_0_2n64sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_2n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_ae34:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "0000";

endmodule

module IFFT_twid_rom_5 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_single_port_rom_5 \gen_auto:rom_component (
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_4(q_a_4),
	.q_a_5(q_a_5),
	.q_a_6(q_a_6),
	.q_a_7(q_a_7),
	.global_clock_enable(global_clock_enable),
	.twad_tdl_0_6(twad_tdl_0_6),
	.twad_tdl_1_6(twad_tdl_1_6),
	.twad_tdl_2_6(twad_tdl_2_6),
	.twad_tdl_3_6(twad_tdl_3_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_single_port_rom_5 (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_4,
	q_a_5,
	q_a_6,
	q_a_7,
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_4;
output 	q_a_5;
output 	q_a_6;
output 	q_a_7;
input 	global_clock_enable;
input 	twad_tdl_0_6;
input 	twad_tdl_1_6;
input 	twad_tdl_2_6;
input 	twad_tdl_3_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_6 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(global_clock_enable),
	.address_a({twad_tdl_3_6,twad_tdl_2_6,twad_tdl_1_6,twad_tdl_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_6 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_be34 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_be34 (
	q_a,
	clocken0,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
input 	clocken0;
input 	[3:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "rom";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "3456";

cyclonev_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "rom";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "F12C";

cyclonev_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "rom";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FA76";

cyclonev_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "rom";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "3760";

cyclonev_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "rom";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "4FF0";

cyclonev_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "rom";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "2AFA";

cyclonev_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "rom";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "19FC";

cyclonev_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain(1'b0),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "IFFT_fft_ii_0_3n64sin.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_3dp_rom:twrom|twid_rom:\\gen_M4K:sin_3n|altera_fft_single_port_rom:\\gen_auto:rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_be34:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "rom";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "F800";

endmodule

module IFFT_asj_fft_4dp_ram (
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_3,
	rdaddress_c_bus_14,
	rdaddress_c_bus_15,
	rdaddress_c_bus_11,
	rdaddress_c_bus_7,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_5,
	ram_in_reg_2_6,
	ram_in_reg_3_3,
	ram_in_reg_3_0,
	ram_in_reg_3_1,
	ram_in_reg_3_2,
	ram_in_reg_3_7,
	ram_in_reg_3_4,
	ram_in_reg_3_5,
	ram_in_reg_3_6,
	ram_in_reg_4_3,
	ram_in_reg_4_0,
	ram_in_reg_4_1,
	ram_in_reg_4_2,
	ram_in_reg_4_7,
	ram_in_reg_4_4,
	ram_in_reg_4_5,
	ram_in_reg_4_6,
	ram_in_reg_5_3,
	ram_in_reg_5_0,
	ram_in_reg_5_1,
	ram_in_reg_5_2,
	ram_in_reg_5_7,
	ram_in_reg_5_4,
	ram_in_reg_5_5,
	ram_in_reg_5_6,
	ram_in_reg_6_3,
	ram_in_reg_6_0,
	ram_in_reg_6_1,
	ram_in_reg_6_2,
	ram_in_reg_6_7,
	ram_in_reg_6_4,
	ram_in_reg_6_5,
	ram_in_reg_6_6,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_1,
	ram_in_reg_7_2,
	ram_in_reg_7_7,
	ram_in_reg_7_4,
	ram_in_reg_7_5,
	ram_in_reg_7_6,
	ram_in_reg_1_31,
	ram_in_reg_1_01,
	ram_in_reg_1_11,
	ram_in_reg_1_21,
	ram_in_reg_1_7,
	ram_in_reg_1_4,
	ram_in_reg_1_5,
	ram_in_reg_1_6,
	ram_in_reg_0_3,
	ram_in_reg_0_01,
	ram_in_reg_0_11,
	ram_in_reg_0_2,
	ram_in_reg_0_7,
	ram_in_reg_0_4,
	ram_in_reg_0_5,
	ram_in_reg_0_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_13;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_3;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_7;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_1;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_7;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_7;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_7;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_7;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_6;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_11;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_asj_fft_data_ram \gen_rams:0:dat_A (
	.q_b_10(q_b_101),
	.q_b_2(q_b_21),
	.q_b_11(q_b_111),
	.q_b_3(q_b_31),
	.q_b_12(q_b_121),
	.q_b_4(q_b_41),
	.q_b_13(q_b_131),
	.q_b_5(q_b_51),
	.q_b_14(q_b_141),
	.q_b_6(q_b_61),
	.q_b_15(q_b_151),
	.q_b_7(q_b_71),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.q_b_9(q_b_91),
	.q_b_1(q_b_16),
	.q_b_8(q_b_81),
	.q_b_0(q_b_01),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_1_01(ram_in_reg_1_01),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_01(ram_in_reg_0_01),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.clk(clk));

IFFT_asj_fft_data_ram_1 \gen_rams:1:dat_A (
	.q_b_10(q_b_102),
	.q_b_2(q_b_22),
	.q_b_11(q_b_112),
	.q_b_3(q_b_32),
	.q_b_12(q_b_122),
	.q_b_4(q_b_42),
	.q_b_13(q_b_132),
	.q_b_5(q_b_52),
	.q_b_14(q_b_142),
	.q_b_6(q_b_62),
	.q_b_15(q_b_152),
	.q_b_7(q_b_72),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.q_b_9(q_b_92),
	.q_b_1(q_b_17),
	.q_b_8(q_b_82),
	.q_b_0(q_b_02),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_1_11(ram_in_reg_1_11),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_11(ram_in_reg_0_11),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.clk(clk));

IFFT_asj_fft_data_ram_3 \gen_rams:3:dat_A (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_3(rdaddress_c_bus_3),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_1_31(ram_in_reg_1_31),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.clk(clk));

IFFT_asj_fft_data_ram_2 \gen_rams:2:dat_A (
	.q_b_10(q_b_103),
	.q_b_2(q_b_23),
	.q_b_11(q_b_113),
	.q_b_3(q_b_33),
	.q_b_12(q_b_123),
	.q_b_4(q_b_43),
	.q_b_13(q_b_133),
	.q_b_5(q_b_53),
	.q_b_14(q_b_143),
	.q_b_6(q_b_63),
	.q_b_15(q_b_153),
	.q_b_7(q_b_73),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_7(rdaddress_c_bus_7),
	.q_b_9(q_b_93),
	.q_b_1(q_b_18),
	.q_b_8(q_b_83),
	.q_b_0(q_b_03),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_1_21(ram_in_reg_1_21),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.clk(clk));

endmodule

module IFFT_asj_fft_data_ram (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_14,
	rdaddress_c_bus_15,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_4,
	ram_in_reg_3_0,
	ram_in_reg_3_4,
	ram_in_reg_4_0,
	ram_in_reg_4_4,
	ram_in_reg_5_0,
	ram_in_reg_5_4,
	ram_in_reg_6_0,
	ram_in_reg_6_4,
	ram_in_reg_7_0,
	ram_in_reg_7_4,
	ram_in_reg_1_01,
	ram_in_reg_1_4,
	ram_in_reg_0_01,
	ram_in_reg_0_4,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_15;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_4;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_4;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_4;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_4;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_1_01(ram_in_reg_1_01),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_01(ram_in_reg_0_01),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_14,
	rdaddress_c_bus_15,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_4,
	ram_in_reg_3_0,
	ram_in_reg_3_4,
	ram_in_reg_4_0,
	ram_in_reg_4_4,
	ram_in_reg_5_0,
	ram_in_reg_5_4,
	ram_in_reg_6_0,
	ram_in_reg_6_4,
	ram_in_reg_7_0,
	ram_in_reg_7_4,
	ram_in_reg_1_01,
	ram_in_reg_1_4,
	ram_in_reg_0_01,
	ram_in_reg_0_4,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_15;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_4;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_4;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_4;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_4;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_7 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wc_vec_3),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_0,ram_in_reg_0_0}),
	.address_b({rdaddress_c_bus_15,rdaddress_c_bus_14,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_0,ram_in_reg_6_0,ram_in_reg_5_0,ram_in_reg_4_0,ram_in_reg_3_0,ram_in_reg_2_0,ram_in_reg_1_01,ram_in_reg_0_01,ram_in_reg_7_4,ram_in_reg_6_4,ram_in_reg_5_4,ram_in_reg_4_4,ram_in_reg_3_4,ram_in_reg_2_4,ram_in_reg_1_4,ram_in_reg_0_4}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_7 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_1 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_5,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_1_11,
	ram_in_reg_1_5,
	ram_in_reg_0_11,
	ram_in_reg_0_5,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_5;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_5;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_11;
input 	ram_in_reg_0_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_1 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_1_11(ram_in_reg_1_11),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_11(ram_in_reg_0_11),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_1 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_11,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_5,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_1_11,
	ram_in_reg_1_5,
	ram_in_reg_0_11,
	ram_in_reg_0_5,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_11;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_5;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_5;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_11;
input 	ram_in_reg_0_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_8 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wc_vec_3),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_1,ram_in_reg_0_1}),
	.address_b({rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_1,ram_in_reg_6_1,ram_in_reg_5_1,ram_in_reg_4_1,ram_in_reg_3_1,ram_in_reg_2_1,ram_in_reg_1_11,ram_in_reg_0_11,ram_in_reg_7_5,ram_in_reg_6_5,ram_in_reg_5_5,ram_in_reg_4_5,ram_in_reg_3_5,ram_in_reg_2_5,ram_in_reg_1_5,ram_in_reg_0_5}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_8 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_1 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_1 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_2 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_14,
	rdaddress_c_bus_7,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_6,
	ram_in_reg_3_2,
	ram_in_reg_3_6,
	ram_in_reg_4_2,
	ram_in_reg_4_6,
	ram_in_reg_5_2,
	ram_in_reg_5_6,
	ram_in_reg_6_2,
	ram_in_reg_6_6,
	ram_in_reg_7_2,
	ram_in_reg_7_6,
	ram_in_reg_1_21,
	ram_in_reg_1_6,
	ram_in_reg_0_2,
	ram_in_reg_0_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_7;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_6;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_2 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_7(rdaddress_c_bus_7),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_1_21(ram_in_reg_1_21),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_2 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_14,
	rdaddress_c_bus_7,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_6,
	ram_in_reg_3_2,
	ram_in_reg_3_6,
	ram_in_reg_4_2,
	ram_in_reg_4_6,
	ram_in_reg_5_2,
	ram_in_reg_5_6,
	ram_in_reg_6_2,
	ram_in_reg_6_6,
	ram_in_reg_7_2,
	ram_in_reg_7_6,
	ram_in_reg_1_21,
	ram_in_reg_1_6,
	ram_in_reg_0_2,
	ram_in_reg_0_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_7;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_6;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_9 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wc_vec_3),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_2,ram_in_reg_0_0}),
	.address_b({rdaddress_c_bus_7,rdaddress_c_bus_14,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_2,ram_in_reg_6_2,ram_in_reg_5_2,ram_in_reg_4_2,ram_in_reg_3_2,ram_in_reg_2_2,ram_in_reg_1_21,ram_in_reg_0_2,ram_in_reg_7_6,ram_in_reg_6_6,ram_in_reg_5_6,ram_in_reg_4_6,ram_in_reg_3_6,ram_in_reg_2_6,ram_in_reg_1_6,ram_in_reg_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_9 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_2 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_2 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_3 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_3,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_7,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_1_31,
	ram_in_reg_1_7,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_3;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_7;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_7;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_7;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_7;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_7;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_7;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_3 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.wc_vec_3(wc_vec_3),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_3(rdaddress_c_bus_3),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_1_31(ram_in_reg_1_31),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_3 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	wc_vec_3,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_3,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_7,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_1_31,
	ram_in_reg_1_7,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	wc_vec_3;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_3;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_7;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_7;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_7;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_7;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_7;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_7;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_10 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wc_vec_3),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_3,ram_in_reg_0_1}),
	.address_b({rdaddress_c_bus_3,rdaddress_c_bus_10,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_3,ram_in_reg_6_3,ram_in_reg_5_3,ram_in_reg_4_3,ram_in_reg_3_3,ram_in_reg_2_3,ram_in_reg_1_31,ram_in_reg_0_3,ram_in_reg_7_7,ram_in_reg_6_7,ram_in_reg_5_7,ram_in_reg_4_7,ram_in_reg_3_7,ram_in_reg_2_7,ram_in_reg_1_7,ram_in_reg_0_7}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_10 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_3 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_3 (
	q_b,
	wren_a,
	address_a,
	address_b,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_C|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_4dp_ram_1 (
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_3,
	wd_vec_3,
	rdaddress_c_bus_14,
	rdaddress_c_bus_15,
	rdaddress_c_bus_11,
	rdaddress_c_bus_7,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_5,
	ram_in_reg_2_6,
	ram_in_reg_3_3,
	ram_in_reg_3_0,
	ram_in_reg_3_1,
	ram_in_reg_3_2,
	ram_in_reg_3_7,
	ram_in_reg_3_4,
	ram_in_reg_3_5,
	ram_in_reg_3_6,
	ram_in_reg_4_3,
	ram_in_reg_4_0,
	ram_in_reg_4_1,
	ram_in_reg_4_2,
	ram_in_reg_4_7,
	ram_in_reg_4_4,
	ram_in_reg_4_5,
	ram_in_reg_4_6,
	ram_in_reg_5_3,
	ram_in_reg_5_0,
	ram_in_reg_5_1,
	ram_in_reg_5_2,
	ram_in_reg_5_7,
	ram_in_reg_5_4,
	ram_in_reg_5_5,
	ram_in_reg_5_6,
	ram_in_reg_6_3,
	ram_in_reg_6_0,
	ram_in_reg_6_1,
	ram_in_reg_6_2,
	ram_in_reg_6_7,
	ram_in_reg_6_4,
	ram_in_reg_6_5,
	ram_in_reg_6_6,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_1,
	ram_in_reg_7_2,
	ram_in_reg_7_7,
	ram_in_reg_7_4,
	ram_in_reg_7_5,
	ram_in_reg_7_6,
	ram_in_reg_1_31,
	ram_in_reg_1_01,
	ram_in_reg_1_11,
	ram_in_reg_1_21,
	ram_in_reg_1_7,
	ram_in_reg_1_4,
	ram_in_reg_1_5,
	ram_in_reg_1_6,
	ram_in_reg_0_3,
	ram_in_reg_0_01,
	ram_in_reg_0_11,
	ram_in_reg_0_2,
	ram_in_reg_0_7,
	ram_in_reg_0_4,
	ram_in_reg_0_5,
	ram_in_reg_0_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_13;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_3;
input 	wd_vec_3;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_15;
input 	rdaddress_c_bus_11;
input 	rdaddress_c_bus_7;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_1;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_7;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_7;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_7;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_7;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_6;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_11;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_asj_fft_data_ram_7 \gen_rams:3:dat_A (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_3(rdaddress_c_bus_3),
	.wd_vec_3(wd_vec_3),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_1_31(ram_in_reg_1_31),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.clk(clk));

IFFT_asj_fft_data_ram_4 \gen_rams:0:dat_A (
	.q_b_10(q_b_101),
	.q_b_2(q_b_21),
	.q_b_11(q_b_111),
	.q_b_3(q_b_31),
	.q_b_12(q_b_121),
	.q_b_4(q_b_41),
	.q_b_13(q_b_131),
	.q_b_5(q_b_51),
	.q_b_14(q_b_141),
	.q_b_6(q_b_61),
	.q_b_15(q_b_151),
	.q_b_7(q_b_71),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.wd_vec_3(wd_vec_3),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.q_b_9(q_b_91),
	.q_b_1(q_b_16),
	.q_b_8(q_b_81),
	.q_b_0(q_b_01),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_1_01(ram_in_reg_1_01),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_01(ram_in_reg_0_01),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.clk(clk));

IFFT_asj_fft_data_ram_5 \gen_rams:1:dat_A (
	.q_b_10(q_b_102),
	.q_b_2(q_b_22),
	.q_b_11(q_b_112),
	.q_b_3(q_b_32),
	.q_b_12(q_b_122),
	.q_b_4(q_b_42),
	.q_b_13(q_b_132),
	.q_b_5(q_b_52),
	.q_b_14(q_b_142),
	.q_b_6(q_b_62),
	.q_b_15(q_b_152),
	.q_b_7(q_b_72),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.wd_vec_3(wd_vec_3),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.q_b_9(q_b_92),
	.q_b_1(q_b_17),
	.q_b_8(q_b_82),
	.q_b_0(q_b_02),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_1_11(ram_in_reg_1_11),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_11(ram_in_reg_0_11),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.clk(clk));

IFFT_asj_fft_data_ram_6 \gen_rams:2:dat_A (
	.q_b_10(q_b_103),
	.q_b_2(q_b_23),
	.q_b_11(q_b_113),
	.q_b_3(q_b_33),
	.q_b_12(q_b_123),
	.q_b_4(q_b_43),
	.q_b_13(q_b_133),
	.q_b_5(q_b_53),
	.q_b_14(q_b_143),
	.q_b_6(q_b_63),
	.q_b_15(q_b_153),
	.q_b_7(q_b_73),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.wd_vec_3(wd_vec_3),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_7(rdaddress_c_bus_7),
	.q_b_9(q_b_93),
	.q_b_1(q_b_18),
	.q_b_8(q_b_83),
	.q_b_0(q_b_03),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_1_21(ram_in_reg_1_21),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.clk(clk));

endmodule

module IFFT_asj_fft_data_ram_4 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	wd_vec_3,
	rdaddress_c_bus_14,
	rdaddress_c_bus_15,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_4,
	ram_in_reg_3_0,
	ram_in_reg_3_4,
	ram_in_reg_4_0,
	ram_in_reg_4_4,
	ram_in_reg_5_0,
	ram_in_reg_5_4,
	ram_in_reg_6_0,
	ram_in_reg_6_4,
	ram_in_reg_7_0,
	ram_in_reg_7_4,
	ram_in_reg_1_01,
	ram_in_reg_1_4,
	ram_in_reg_0_01,
	ram_in_reg_0_4,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	wd_vec_3;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_15;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_4;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_4;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_4;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_4;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_4 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.wd_vec_3(wd_vec_3),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_15(rdaddress_c_bus_15),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_1_01(ram_in_reg_1_01),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.ram_in_reg_0_01(ram_in_reg_0_01),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_4 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	wd_vec_3,
	rdaddress_c_bus_14,
	rdaddress_c_bus_15,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_4,
	ram_in_reg_3_0,
	ram_in_reg_3_4,
	ram_in_reg_4_0,
	ram_in_reg_4_4,
	ram_in_reg_5_0,
	ram_in_reg_5_4,
	ram_in_reg_6_0,
	ram_in_reg_6_4,
	ram_in_reg_7_0,
	ram_in_reg_7_4,
	ram_in_reg_1_01,
	ram_in_reg_1_4,
	ram_in_reg_0_01,
	ram_in_reg_0_4,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	wd_vec_3;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_15;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_4;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_4;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_4;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_4;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_4;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_4;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_11 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_0,ram_in_reg_0_0}),
	.address_b({rdaddress_c_bus_15,rdaddress_c_bus_14,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.wren_a(wd_vec_3),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_0,ram_in_reg_6_0,ram_in_reg_5_0,ram_in_reg_4_0,ram_in_reg_3_0,ram_in_reg_2_0,ram_in_reg_1_01,ram_in_reg_0_01,ram_in_reg_7_4,ram_in_reg_6_4,ram_in_reg_5_4,ram_in_reg_4_4,ram_in_reg_3_4,ram_in_reg_2_4,ram_in_reg_1_4,ram_in_reg_0_4}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_11 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_4 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_4 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_5 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	wd_vec_3,
	rdaddress_c_bus_11,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_5,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_1_11,
	ram_in_reg_1_5,
	ram_in_reg_0_11,
	ram_in_reg_0_5,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	wd_vec_3;
input 	rdaddress_c_bus_11;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_5;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_5;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_11;
input 	ram_in_reg_0_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_5 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.wd_vec_3(wd_vec_3),
	.rdaddress_c_bus_11(rdaddress_c_bus_11),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_1_11(ram_in_reg_1_11),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_11(ram_in_reg_0_11),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_5 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	wd_vec_3,
	rdaddress_c_bus_11,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_5,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_1_11,
	ram_in_reg_1_5,
	ram_in_reg_0_11,
	ram_in_reg_0_5,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	wd_vec_3;
input 	rdaddress_c_bus_11;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_5;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_5;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_11;
input 	ram_in_reg_0_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_12 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_1,ram_in_reg_0_1}),
	.address_b({rdaddress_c_bus_11,rdaddress_c_bus_10,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.wren_a(wd_vec_3),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_1,ram_in_reg_6_1,ram_in_reg_5_1,ram_in_reg_4_1,ram_in_reg_3_1,ram_in_reg_2_1,ram_in_reg_1_11,ram_in_reg_0_11,ram_in_reg_7_5,ram_in_reg_6_5,ram_in_reg_5_5,ram_in_reg_4_5,ram_in_reg_3_5,ram_in_reg_2_5,ram_in_reg_1_5,ram_in_reg_0_5}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_12 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_5 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_5 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_6 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	wd_vec_3,
	rdaddress_c_bus_14,
	rdaddress_c_bus_7,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_6,
	ram_in_reg_3_2,
	ram_in_reg_3_6,
	ram_in_reg_4_2,
	ram_in_reg_4_6,
	ram_in_reg_5_2,
	ram_in_reg_5_6,
	ram_in_reg_6_2,
	ram_in_reg_6_6,
	ram_in_reg_7_2,
	ram_in_reg_7_6,
	ram_in_reg_1_21,
	ram_in_reg_1_6,
	ram_in_reg_0_2,
	ram_in_reg_0_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	wd_vec_3;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_7;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_6;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_6 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.wd_vec_3(wd_vec_3),
	.rdaddress_c_bus_14(rdaddress_c_bus_14),
	.rdaddress_c_bus_7(rdaddress_c_bus_7),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_1_21(ram_in_reg_1_21),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_6 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	wd_vec_3,
	rdaddress_c_bus_14,
	rdaddress_c_bus_7,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_6,
	ram_in_reg_3_2,
	ram_in_reg_3_6,
	ram_in_reg_4_2,
	ram_in_reg_4_6,
	ram_in_reg_5_2,
	ram_in_reg_5_6,
	ram_in_reg_6_2,
	ram_in_reg_6_6,
	ram_in_reg_7_2,
	ram_in_reg_7_6,
	ram_in_reg_1_21,
	ram_in_reg_1_6,
	ram_in_reg_0_2,
	ram_in_reg_0_6,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	wd_vec_3;
input 	rdaddress_c_bus_14;
input 	rdaddress_c_bus_7;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_0_0;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_6;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_13 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_2,ram_in_reg_0_0}),
	.address_b({rdaddress_c_bus_7,rdaddress_c_bus_14,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.wren_a(wd_vec_3),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_2,ram_in_reg_6_2,ram_in_reg_5_2,ram_in_reg_4_2,ram_in_reg_3_2,ram_in_reg_2_2,ram_in_reg_1_21,ram_in_reg_0_2,ram_in_reg_7_6,ram_in_reg_6_6,ram_in_reg_5_6,ram_in_reg_4_6,ram_in_reg_3_6,ram_in_reg_2_6,ram_in_reg_1_6,ram_in_reg_0_6}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_13 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_6 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_6 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_7 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_3,
	wd_vec_3,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_7,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_1_31,
	ram_in_reg_1_7,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_3;
input 	wd_vec_3;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_7;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_7;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_7;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_7;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_7;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_7;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_7 \gen_M4K:ram_component (
	.q_b_10(q_b_10),
	.q_b_2(q_b_2),
	.q_b_11(q_b_11),
	.q_b_3(q_b_3),
	.q_b_12(q_b_12),
	.q_b_4(q_b_4),
	.q_b_13(q_b_13),
	.q_b_5(q_b_5),
	.q_b_14(q_b_14),
	.q_b_6(q_b_6),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.ram_block6a0(ram_block6a0),
	.ram_block6a1(ram_block6a1),
	.rdaddress_c_bus_0(rdaddress_c_bus_0),
	.rdaddress_c_bus_13(rdaddress_c_bus_13),
	.rdaddress_c_bus_10(rdaddress_c_bus_10),
	.rdaddress_c_bus_3(rdaddress_c_bus_3),
	.wd_vec_3(wd_vec_3),
	.q_b_9(q_b_9),
	.q_b_1(q_b_1),
	.q_b_8(q_b_8),
	.q_b_0(q_b_0),
	.global_clock_enable(global_clock_enable),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_1_31(ram_in_reg_1_31),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_7 (
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_13,
	q_b_5,
	q_b_14,
	q_b_6,
	q_b_15,
	q_b_7,
	ram_block6a0,
	ram_block6a1,
	rdaddress_c_bus_0,
	rdaddress_c_bus_13,
	rdaddress_c_bus_10,
	rdaddress_c_bus_3,
	wd_vec_3,
	q_b_9,
	q_b_1,
	q_b_8,
	q_b_0,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_7,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_1_31,
	ram_in_reg_1_7,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_13;
output 	q_b_5;
output 	q_b_14;
output 	q_b_6;
output 	q_b_15;
output 	q_b_7;
input 	ram_block6a0;
input 	ram_block6a1;
input 	rdaddress_c_bus_0;
input 	rdaddress_c_bus_13;
input 	rdaddress_c_bus_10;
input 	rdaddress_c_bus_3;
input 	wd_vec_3;
output 	q_b_9;
output 	q_b_1;
output 	q_b_8;
output 	q_b_0;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_7;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_7;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_7;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_7;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_7;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_7;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_7;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_14 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({ram_block6a1,ram_block6a0,ram_in_reg_1_3,ram_in_reg_0_1}),
	.address_b({rdaddress_c_bus_3,rdaddress_c_bus_10,rdaddress_c_bus_13,rdaddress_c_bus_0}),
	.wren_a(wd_vec_3),
	.clocken0(global_clock_enable),
	.data_a({ram_in_reg_7_3,ram_in_reg_6_3,ram_in_reg_5_3,ram_in_reg_4_3,ram_in_reg_3_3,ram_in_reg_2_3,ram_in_reg_1_31,ram_in_reg_0_3,ram_in_reg_7_7,ram_in_reg_6_7,ram_in_reg_5_7,ram_in_reg_4_7,ram_in_reg_3_7,ram_in_reg_2_7,ram_in_reg_1_7,ram_in_reg_0_7}),
	.clock0(clk));

endmodule

module IFFT_altsyncram_14 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_7 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_7 (
	q_b,
	address_a,
	address_b,
	wren_a,
	clocken0,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	clocken0;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:\\gen_M4K_Output:dat_D|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_4dp_ram_2 (
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	wren_a_1,
	a_ram_data_in_bus_46,
	wraddress_a_bus_0,
	wraddress_a_bus_9,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_0,
	rdaddress_a_bus_9,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wren_a_2,
	a_ram_data_in_bus_30,
	wraddress_a_bus_12,
	wraddress_a_bus_5,
	rdaddress_a_bus_12,
	rdaddress_a_bus_5,
	wren_a_3,
	a_ram_data_in_bus_14,
	wraddress_a_bus_1,
	rdaddress_a_bus_1,
	wren_a_0,
	a_ram_data_in_bus_62,
	wraddress_a_bus_13,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_52,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_32,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_1,
	a_ram_data_in_bus_49,
	a_ram_data_in_bus_33,
	a_ram_data_in_bus_17,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_13;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
output 	q_b_1;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
input 	wren_a_1;
input 	a_ram_data_in_bus_46;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_9;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_9;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wren_a_2;
input 	a_ram_data_in_bus_30;
input 	wraddress_a_bus_12;
input 	wraddress_a_bus_5;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_5;
input 	wren_a_3;
input 	a_ram_data_in_bus_14;
input 	wraddress_a_bus_1;
input 	rdaddress_a_bus_1;
input 	wren_a_0;
input 	a_ram_data_in_bus_62;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_42;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_58;
input 	a_ram_data_in_bus_43;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_63;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_52;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_0;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_32;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_1;
input 	a_ram_data_in_bus_49;
input 	a_ram_data_in_bus_33;
input 	a_ram_data_in_bus_17;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_asj_fft_data_ram_8 \gen_rams:0:dat_A (
	.q_b_14(q_b_143),
	.q_b_13(q_b_133),
	.q_b_10(q_b_103),
	.q_b_11(q_b_113),
	.q_b_12(q_b_123),
	.q_b_15(q_b_153),
	.q_b_7(q_b_73),
	.q_b_6(q_b_63),
	.q_b_3(q_b_33),
	.q_b_4(q_b_43),
	.q_b_5(q_b_53),
	.q_b_2(q_b_23),
	.q_b_8(q_b_82),
	.q_b_9(q_b_92),
	.q_b_0(q_b_01),
	.q_b_1(q_b_16),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.wren_a_0(wren_a_0),
	.a_ram_data_in_bus_62(a_ram_data_in_bus_62),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.a_ram_data_in_bus_61(a_ram_data_in_bus_61),
	.a_ram_data_in_bus_58(a_ram_data_in_bus_58),
	.a_ram_data_in_bus_59(a_ram_data_in_bus_59),
	.a_ram_data_in_bus_60(a_ram_data_in_bus_60),
	.a_ram_data_in_bus_63(a_ram_data_in_bus_63),
	.a_ram_data_in_bus_55(a_ram_data_in_bus_55),
	.a_ram_data_in_bus_54(a_ram_data_in_bus_54),
	.a_ram_data_in_bus_51(a_ram_data_in_bus_51),
	.a_ram_data_in_bus_52(a_ram_data_in_bus_52),
	.a_ram_data_in_bus_53(a_ram_data_in_bus_53),
	.a_ram_data_in_bus_50(a_ram_data_in_bus_50),
	.a_ram_data_in_bus_56(a_ram_data_in_bus_56),
	.a_ram_data_in_bus_57(a_ram_data_in_bus_57),
	.a_ram_data_in_bus_48(a_ram_data_in_bus_48),
	.a_ram_data_in_bus_49(a_ram_data_in_bus_49),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

IFFT_asj_fft_data_ram_9 \gen_rams:1:dat_A (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_83),
	.q_b_9(q_b_93),
	.q_b_0(q_b_02),
	.q_b_1(q_b_17),
	.wren_a_1(wren_a_1),
	.a_ram_data_in_bus_46(a_ram_data_in_bus_46),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_9(wraddress_a_bus_9),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_9(rdaddress_a_bus_9),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.a_ram_data_in_bus_45(a_ram_data_in_bus_45),
	.a_ram_data_in_bus_42(a_ram_data_in_bus_42),
	.a_ram_data_in_bus_43(a_ram_data_in_bus_43),
	.a_ram_data_in_bus_44(a_ram_data_in_bus_44),
	.a_ram_data_in_bus_47(a_ram_data_in_bus_47),
	.a_ram_data_in_bus_39(a_ram_data_in_bus_39),
	.a_ram_data_in_bus_38(a_ram_data_in_bus_38),
	.a_ram_data_in_bus_35(a_ram_data_in_bus_35),
	.a_ram_data_in_bus_36(a_ram_data_in_bus_36),
	.a_ram_data_in_bus_37(a_ram_data_in_bus_37),
	.a_ram_data_in_bus_34(a_ram_data_in_bus_34),
	.a_ram_data_in_bus_40(a_ram_data_in_bus_40),
	.a_ram_data_in_bus_41(a_ram_data_in_bus_41),
	.a_ram_data_in_bus_32(a_ram_data_in_bus_32),
	.a_ram_data_in_bus_33(a_ram_data_in_bus_33),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

IFFT_asj_fft_data_ram_11 \gen_rams:3:dat_A (
	.q_b_14(q_b_142),
	.q_b_13(q_b_132),
	.q_b_10(q_b_102),
	.q_b_11(q_b_112),
	.q_b_12(q_b_122),
	.q_b_15(q_b_152),
	.q_b_7(q_b_72),
	.q_b_6(q_b_62),
	.q_b_3(q_b_32),
	.q_b_4(q_b_42),
	.q_b_5(q_b_52),
	.q_b_2(q_b_22),
	.q_b_8(q_b_81),
	.q_b_9(q_b_91),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.wren_a_3(wren_a_3),
	.a_ram_data_in_bus_14(a_ram_data_in_bus_14),
	.wraddress_a_bus_1(wraddress_a_bus_1),
	.rdaddress_a_bus_1(rdaddress_a_bus_1),
	.a_ram_data_in_bus_13(a_ram_data_in_bus_13),
	.a_ram_data_in_bus_10(a_ram_data_in_bus_10),
	.a_ram_data_in_bus_11(a_ram_data_in_bus_11),
	.a_ram_data_in_bus_12(a_ram_data_in_bus_12),
	.a_ram_data_in_bus_15(a_ram_data_in_bus_15),
	.a_ram_data_in_bus_7(a_ram_data_in_bus_7),
	.a_ram_data_in_bus_6(a_ram_data_in_bus_6),
	.a_ram_data_in_bus_3(a_ram_data_in_bus_3),
	.a_ram_data_in_bus_4(a_ram_data_in_bus_4),
	.a_ram_data_in_bus_5(a_ram_data_in_bus_5),
	.a_ram_data_in_bus_2(a_ram_data_in_bus_2),
	.a_ram_data_in_bus_8(a_ram_data_in_bus_8),
	.a_ram_data_in_bus_9(a_ram_data_in_bus_9),
	.a_ram_data_in_bus_0(a_ram_data_in_bus_0),
	.a_ram_data_in_bus_1(a_ram_data_in_bus_1),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

IFFT_asj_fft_data_ram_10 \gen_rams:2:dat_A (
	.q_b_14(q_b_141),
	.q_b_13(q_b_131),
	.q_b_10(q_b_101),
	.q_b_11(q_b_111),
	.q_b_12(q_b_121),
	.q_b_15(q_b_151),
	.q_b_7(q_b_71),
	.q_b_6(q_b_61),
	.q_b_3(q_b_31),
	.q_b_4(q_b_41),
	.q_b_5(q_b_51),
	.q_b_2(q_b_21),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_03),
	.q_b_1(q_b_18),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.wren_a_2(wren_a_2),
	.a_ram_data_in_bus_30(a_ram_data_in_bus_30),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.wraddress_a_bus_5(wraddress_a_bus_5),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.rdaddress_a_bus_5(rdaddress_a_bus_5),
	.a_ram_data_in_bus_29(a_ram_data_in_bus_29),
	.a_ram_data_in_bus_26(a_ram_data_in_bus_26),
	.a_ram_data_in_bus_27(a_ram_data_in_bus_27),
	.a_ram_data_in_bus_28(a_ram_data_in_bus_28),
	.a_ram_data_in_bus_31(a_ram_data_in_bus_31),
	.a_ram_data_in_bus_23(a_ram_data_in_bus_23),
	.a_ram_data_in_bus_22(a_ram_data_in_bus_22),
	.a_ram_data_in_bus_19(a_ram_data_in_bus_19),
	.a_ram_data_in_bus_20(a_ram_data_in_bus_20),
	.a_ram_data_in_bus_21(a_ram_data_in_bus_21),
	.a_ram_data_in_bus_18(a_ram_data_in_bus_18),
	.a_ram_data_in_bus_24(a_ram_data_in_bus_24),
	.a_ram_data_in_bus_25(a_ram_data_in_bus_25),
	.a_ram_data_in_bus_16(a_ram_data_in_bus_16),
	.a_ram_data_in_bus_17(a_ram_data_in_bus_17),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_asj_fft_data_ram_8 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wraddress_a_bus_12,
	rdaddress_a_bus_12,
	wren_a_0,
	a_ram_data_in_bus_62,
	wraddress_a_bus_13,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_52,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_49,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wraddress_a_bus_12;
input 	rdaddress_a_bus_12;
input 	wren_a_0;
input 	a_ram_data_in_bus_62;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_58;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_63;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_52;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_49;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_8 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.wren_a_0(wren_a_0),
	.a_ram_data_in_bus_62(a_ram_data_in_bus_62),
	.wraddress_a_bus_13(wraddress_a_bus_13),
	.rdaddress_a_bus_13(rdaddress_a_bus_13),
	.a_ram_data_in_bus_61(a_ram_data_in_bus_61),
	.a_ram_data_in_bus_58(a_ram_data_in_bus_58),
	.a_ram_data_in_bus_59(a_ram_data_in_bus_59),
	.a_ram_data_in_bus_60(a_ram_data_in_bus_60),
	.a_ram_data_in_bus_63(a_ram_data_in_bus_63),
	.a_ram_data_in_bus_55(a_ram_data_in_bus_55),
	.a_ram_data_in_bus_54(a_ram_data_in_bus_54),
	.a_ram_data_in_bus_51(a_ram_data_in_bus_51),
	.a_ram_data_in_bus_52(a_ram_data_in_bus_52),
	.a_ram_data_in_bus_53(a_ram_data_in_bus_53),
	.a_ram_data_in_bus_50(a_ram_data_in_bus_50),
	.a_ram_data_in_bus_56(a_ram_data_in_bus_56),
	.a_ram_data_in_bus_57(a_ram_data_in_bus_57),
	.a_ram_data_in_bus_48(a_ram_data_in_bus_48),
	.a_ram_data_in_bus_49(a_ram_data_in_bus_49),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_8 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wraddress_a_bus_12,
	rdaddress_a_bus_12,
	wren_a_0,
	a_ram_data_in_bus_62,
	wraddress_a_bus_13,
	rdaddress_a_bus_13,
	a_ram_data_in_bus_61,
	a_ram_data_in_bus_58,
	a_ram_data_in_bus_59,
	a_ram_data_in_bus_60,
	a_ram_data_in_bus_63,
	a_ram_data_in_bus_55,
	a_ram_data_in_bus_54,
	a_ram_data_in_bus_51,
	a_ram_data_in_bus_52,
	a_ram_data_in_bus_53,
	a_ram_data_in_bus_50,
	a_ram_data_in_bus_56,
	a_ram_data_in_bus_57,
	a_ram_data_in_bus_48,
	a_ram_data_in_bus_49,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wraddress_a_bus_12;
input 	rdaddress_a_bus_12;
input 	wren_a_0;
input 	a_ram_data_in_bus_62;
input 	wraddress_a_bus_13;
input 	rdaddress_a_bus_13;
input 	a_ram_data_in_bus_61;
input 	a_ram_data_in_bus_58;
input 	a_ram_data_in_bus_59;
input 	a_ram_data_in_bus_60;
input 	a_ram_data_in_bus_63;
input 	a_ram_data_in_bus_55;
input 	a_ram_data_in_bus_54;
input 	a_ram_data_in_bus_51;
input 	a_ram_data_in_bus_52;
input 	a_ram_data_in_bus_53;
input 	a_ram_data_in_bus_50;
input 	a_ram_data_in_bus_56;
input 	a_ram_data_in_bus_57;
input 	a_ram_data_in_bus_48;
input 	a_ram_data_in_bus_49;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_15 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({wraddress_a_bus_11,wraddress_a_bus_10,wraddress_a_bus_13,wraddress_a_bus_12}),
	.address_b({rdaddress_a_bus_11,rdaddress_a_bus_10,rdaddress_a_bus_13,rdaddress_a_bus_12}),
	.wren_a(wren_a_0),
	.data_a({a_ram_data_in_bus_63,a_ram_data_in_bus_62,a_ram_data_in_bus_61,a_ram_data_in_bus_60,a_ram_data_in_bus_59,a_ram_data_in_bus_58,a_ram_data_in_bus_57,a_ram_data_in_bus_56,a_ram_data_in_bus_55,a_ram_data_in_bus_54,a_ram_data_in_bus_53,a_ram_data_in_bus_52,
a_ram_data_in_bus_51,a_ram_data_in_bus_50,a_ram_data_in_bus_49,a_ram_data_in_bus_48}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_15 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_8 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_8 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_9 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wren_a_1,
	a_ram_data_in_bus_46,
	wraddress_a_bus_0,
	wraddress_a_bus_9,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_0,
	rdaddress_a_bus_9,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_32,
	a_ram_data_in_bus_33,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wren_a_1;
input 	a_ram_data_in_bus_46;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_9;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_9;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_42;
input 	a_ram_data_in_bus_43;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_32;
input 	a_ram_data_in_bus_33;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_9 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wren_a_1(wren_a_1),
	.a_ram_data_in_bus_46(a_ram_data_in_bus_46),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_9(wraddress_a_bus_9),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_9(rdaddress_a_bus_9),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.a_ram_data_in_bus_45(a_ram_data_in_bus_45),
	.a_ram_data_in_bus_42(a_ram_data_in_bus_42),
	.a_ram_data_in_bus_43(a_ram_data_in_bus_43),
	.a_ram_data_in_bus_44(a_ram_data_in_bus_44),
	.a_ram_data_in_bus_47(a_ram_data_in_bus_47),
	.a_ram_data_in_bus_39(a_ram_data_in_bus_39),
	.a_ram_data_in_bus_38(a_ram_data_in_bus_38),
	.a_ram_data_in_bus_35(a_ram_data_in_bus_35),
	.a_ram_data_in_bus_36(a_ram_data_in_bus_36),
	.a_ram_data_in_bus_37(a_ram_data_in_bus_37),
	.a_ram_data_in_bus_34(a_ram_data_in_bus_34),
	.a_ram_data_in_bus_40(a_ram_data_in_bus_40),
	.a_ram_data_in_bus_41(a_ram_data_in_bus_41),
	.a_ram_data_in_bus_32(a_ram_data_in_bus_32),
	.a_ram_data_in_bus_33(a_ram_data_in_bus_33),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_9 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wren_a_1,
	a_ram_data_in_bus_46,
	wraddress_a_bus_0,
	wraddress_a_bus_9,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_0,
	rdaddress_a_bus_9,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	a_ram_data_in_bus_45,
	a_ram_data_in_bus_42,
	a_ram_data_in_bus_43,
	a_ram_data_in_bus_44,
	a_ram_data_in_bus_47,
	a_ram_data_in_bus_39,
	a_ram_data_in_bus_38,
	a_ram_data_in_bus_35,
	a_ram_data_in_bus_36,
	a_ram_data_in_bus_37,
	a_ram_data_in_bus_34,
	a_ram_data_in_bus_40,
	a_ram_data_in_bus_41,
	a_ram_data_in_bus_32,
	a_ram_data_in_bus_33,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wren_a_1;
input 	a_ram_data_in_bus_46;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_9;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_9;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	a_ram_data_in_bus_45;
input 	a_ram_data_in_bus_42;
input 	a_ram_data_in_bus_43;
input 	a_ram_data_in_bus_44;
input 	a_ram_data_in_bus_47;
input 	a_ram_data_in_bus_39;
input 	a_ram_data_in_bus_38;
input 	a_ram_data_in_bus_35;
input 	a_ram_data_in_bus_36;
input 	a_ram_data_in_bus_37;
input 	a_ram_data_in_bus_34;
input 	a_ram_data_in_bus_40;
input 	a_ram_data_in_bus_41;
input 	a_ram_data_in_bus_32;
input 	a_ram_data_in_bus_33;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_16 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_a_1),
	.data_a({a_ram_data_in_bus_47,a_ram_data_in_bus_46,a_ram_data_in_bus_45,a_ram_data_in_bus_44,a_ram_data_in_bus_43,a_ram_data_in_bus_42,a_ram_data_in_bus_41,a_ram_data_in_bus_40,a_ram_data_in_bus_39,a_ram_data_in_bus_38,a_ram_data_in_bus_37,a_ram_data_in_bus_36,
a_ram_data_in_bus_35,a_ram_data_in_bus_34,a_ram_data_in_bus_33,a_ram_data_in_bus_32}),
	.address_a({wraddress_a_bus_11,wraddress_a_bus_10,wraddress_a_bus_9,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_11,rdaddress_a_bus_10,rdaddress_a_bus_9,rdaddress_a_bus_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_16 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[15:0] data_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_9 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_9 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[15:0] data_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_10 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wren_a_2,
	a_ram_data_in_bus_30,
	wraddress_a_bus_12,
	wraddress_a_bus_5,
	rdaddress_a_bus_12,
	rdaddress_a_bus_5,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_17,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wren_a_2;
input 	a_ram_data_in_bus_30;
input 	wraddress_a_bus_12;
input 	wraddress_a_bus_5;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_5;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_17;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_10 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.wren_a_2(wren_a_2),
	.a_ram_data_in_bus_30(a_ram_data_in_bus_30),
	.wraddress_a_bus_12(wraddress_a_bus_12),
	.wraddress_a_bus_5(wraddress_a_bus_5),
	.rdaddress_a_bus_12(rdaddress_a_bus_12),
	.rdaddress_a_bus_5(rdaddress_a_bus_5),
	.a_ram_data_in_bus_29(a_ram_data_in_bus_29),
	.a_ram_data_in_bus_26(a_ram_data_in_bus_26),
	.a_ram_data_in_bus_27(a_ram_data_in_bus_27),
	.a_ram_data_in_bus_28(a_ram_data_in_bus_28),
	.a_ram_data_in_bus_31(a_ram_data_in_bus_31),
	.a_ram_data_in_bus_23(a_ram_data_in_bus_23),
	.a_ram_data_in_bus_22(a_ram_data_in_bus_22),
	.a_ram_data_in_bus_19(a_ram_data_in_bus_19),
	.a_ram_data_in_bus_20(a_ram_data_in_bus_20),
	.a_ram_data_in_bus_21(a_ram_data_in_bus_21),
	.a_ram_data_in_bus_18(a_ram_data_in_bus_18),
	.a_ram_data_in_bus_24(a_ram_data_in_bus_24),
	.a_ram_data_in_bus_25(a_ram_data_in_bus_25),
	.a_ram_data_in_bus_16(a_ram_data_in_bus_16),
	.a_ram_data_in_bus_17(a_ram_data_in_bus_17),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_10 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wren_a_2,
	a_ram_data_in_bus_30,
	wraddress_a_bus_12,
	wraddress_a_bus_5,
	rdaddress_a_bus_12,
	rdaddress_a_bus_5,
	a_ram_data_in_bus_29,
	a_ram_data_in_bus_26,
	a_ram_data_in_bus_27,
	a_ram_data_in_bus_28,
	a_ram_data_in_bus_31,
	a_ram_data_in_bus_23,
	a_ram_data_in_bus_22,
	a_ram_data_in_bus_19,
	a_ram_data_in_bus_20,
	a_ram_data_in_bus_21,
	a_ram_data_in_bus_18,
	a_ram_data_in_bus_24,
	a_ram_data_in_bus_25,
	a_ram_data_in_bus_16,
	a_ram_data_in_bus_17,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wren_a_2;
input 	a_ram_data_in_bus_30;
input 	wraddress_a_bus_12;
input 	wraddress_a_bus_5;
input 	rdaddress_a_bus_12;
input 	rdaddress_a_bus_5;
input 	a_ram_data_in_bus_29;
input 	a_ram_data_in_bus_26;
input 	a_ram_data_in_bus_27;
input 	a_ram_data_in_bus_28;
input 	a_ram_data_in_bus_31;
input 	a_ram_data_in_bus_23;
input 	a_ram_data_in_bus_22;
input 	a_ram_data_in_bus_19;
input 	a_ram_data_in_bus_20;
input 	a_ram_data_in_bus_21;
input 	a_ram_data_in_bus_18;
input 	a_ram_data_in_bus_24;
input 	a_ram_data_in_bus_25;
input 	a_ram_data_in_bus_16;
input 	a_ram_data_in_bus_17;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_17 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({wraddress_a_bus_11,wraddress_a_bus_10,wraddress_a_bus_5,wraddress_a_bus_12}),
	.address_b({rdaddress_a_bus_11,rdaddress_a_bus_10,rdaddress_a_bus_5,rdaddress_a_bus_12}),
	.wren_a(wren_a_2),
	.data_a({a_ram_data_in_bus_31,a_ram_data_in_bus_30,a_ram_data_in_bus_29,a_ram_data_in_bus_28,a_ram_data_in_bus_27,a_ram_data_in_bus_26,a_ram_data_in_bus_25,a_ram_data_in_bus_24,a_ram_data_in_bus_23,a_ram_data_in_bus_22,a_ram_data_in_bus_21,a_ram_data_in_bus_20,
a_ram_data_in_bus_19,a_ram_data_in_bus_18,a_ram_data_in_bus_17,a_ram_data_in_bus_16}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_17 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_10 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_10 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_11 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_a_bus_0,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_0,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wren_a_3,
	a_ram_data_in_bus_14,
	wraddress_a_bus_1,
	rdaddress_a_bus_1,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_1,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wren_a_3;
input 	a_ram_data_in_bus_14;
input 	wraddress_a_bus_1;
input 	rdaddress_a_bus_1;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_0;
input 	a_ram_data_in_bus_1;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_11 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_a_bus_0(wraddress_a_bus_0),
	.wraddress_a_bus_10(wraddress_a_bus_10),
	.wraddress_a_bus_11(wraddress_a_bus_11),
	.rdaddress_a_bus_0(rdaddress_a_bus_0),
	.rdaddress_a_bus_10(rdaddress_a_bus_10),
	.rdaddress_a_bus_11(rdaddress_a_bus_11),
	.wren_a_3(wren_a_3),
	.a_ram_data_in_bus_14(a_ram_data_in_bus_14),
	.wraddress_a_bus_1(wraddress_a_bus_1),
	.rdaddress_a_bus_1(rdaddress_a_bus_1),
	.a_ram_data_in_bus_13(a_ram_data_in_bus_13),
	.a_ram_data_in_bus_10(a_ram_data_in_bus_10),
	.a_ram_data_in_bus_11(a_ram_data_in_bus_11),
	.a_ram_data_in_bus_12(a_ram_data_in_bus_12),
	.a_ram_data_in_bus_15(a_ram_data_in_bus_15),
	.a_ram_data_in_bus_7(a_ram_data_in_bus_7),
	.a_ram_data_in_bus_6(a_ram_data_in_bus_6),
	.a_ram_data_in_bus_3(a_ram_data_in_bus_3),
	.a_ram_data_in_bus_4(a_ram_data_in_bus_4),
	.a_ram_data_in_bus_5(a_ram_data_in_bus_5),
	.a_ram_data_in_bus_2(a_ram_data_in_bus_2),
	.a_ram_data_in_bus_8(a_ram_data_in_bus_8),
	.a_ram_data_in_bus_9(a_ram_data_in_bus_9),
	.a_ram_data_in_bus_0(a_ram_data_in_bus_0),
	.a_ram_data_in_bus_1(a_ram_data_in_bus_1),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_11 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_a_bus_0,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_0,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	wren_a_3,
	a_ram_data_in_bus_14,
	wraddress_a_bus_1,
	rdaddress_a_bus_1,
	a_ram_data_in_bus_13,
	a_ram_data_in_bus_10,
	a_ram_data_in_bus_11,
	a_ram_data_in_bus_12,
	a_ram_data_in_bus_15,
	a_ram_data_in_bus_7,
	a_ram_data_in_bus_6,
	a_ram_data_in_bus_3,
	a_ram_data_in_bus_4,
	a_ram_data_in_bus_5,
	a_ram_data_in_bus_2,
	a_ram_data_in_bus_8,
	a_ram_data_in_bus_9,
	a_ram_data_in_bus_0,
	a_ram_data_in_bus_1,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_a_bus_0;
input 	wraddress_a_bus_10;
input 	wraddress_a_bus_11;
input 	rdaddress_a_bus_0;
input 	rdaddress_a_bus_10;
input 	rdaddress_a_bus_11;
input 	wren_a_3;
input 	a_ram_data_in_bus_14;
input 	wraddress_a_bus_1;
input 	rdaddress_a_bus_1;
input 	a_ram_data_in_bus_13;
input 	a_ram_data_in_bus_10;
input 	a_ram_data_in_bus_11;
input 	a_ram_data_in_bus_12;
input 	a_ram_data_in_bus_15;
input 	a_ram_data_in_bus_7;
input 	a_ram_data_in_bus_6;
input 	a_ram_data_in_bus_3;
input 	a_ram_data_in_bus_4;
input 	a_ram_data_in_bus_5;
input 	a_ram_data_in_bus_2;
input 	a_ram_data_in_bus_8;
input 	a_ram_data_in_bus_9;
input 	a_ram_data_in_bus_0;
input 	a_ram_data_in_bus_1;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_18 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({wraddress_a_bus_11,wraddress_a_bus_10,wraddress_a_bus_1,wraddress_a_bus_0}),
	.address_b({rdaddress_a_bus_11,rdaddress_a_bus_10,rdaddress_a_bus_1,rdaddress_a_bus_0}),
	.wren_a(wren_a_3),
	.data_a({a_ram_data_in_bus_15,a_ram_data_in_bus_14,a_ram_data_in_bus_13,a_ram_data_in_bus_12,a_ram_data_in_bus_11,a_ram_data_in_bus_10,a_ram_data_in_bus_9,a_ram_data_in_bus_8,a_ram_data_in_bus_7,a_ram_data_in_bus_6,a_ram_data_in_bus_5,a_ram_data_in_bus_4,a_ram_data_in_bus_3,
a_ram_data_in_bus_2,a_ram_data_in_bus_1,a_ram_data_in_bus_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_18 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_11 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_11 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_A|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_4dp_ram_3 (
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	wren_b_1,
	b_ram_data_in_bus_46,
	wraddress_b_bus_0,
	wraddress_b_bus_9,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_0,
	rdaddress_b_bus_9,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wren_b_2,
	b_ram_data_in_bus_30,
	wraddress_b_bus_12,
	wraddress_b_bus_5,
	rdaddress_b_bus_12,
	rdaddress_b_bus_5,
	wren_b_3,
	b_ram_data_in_bus_14,
	wraddress_b_bus_1,
	rdaddress_b_bus_1,
	wren_b_0,
	b_ram_data_in_bus_62,
	wraddress_b_bus_13,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_45,
	b_ram_data_in_bus_29,
	b_ram_data_in_bus_13,
	b_ram_data_in_bus_61,
	b_ram_data_in_bus_42,
	b_ram_data_in_bus_26,
	b_ram_data_in_bus_10,
	b_ram_data_in_bus_58,
	b_ram_data_in_bus_43,
	b_ram_data_in_bus_27,
	b_ram_data_in_bus_11,
	b_ram_data_in_bus_59,
	b_ram_data_in_bus_44,
	b_ram_data_in_bus_28,
	b_ram_data_in_bus_12,
	b_ram_data_in_bus_60,
	b_ram_data_in_bus_47,
	b_ram_data_in_bus_31,
	b_ram_data_in_bus_15,
	b_ram_data_in_bus_63,
	b_ram_data_in_bus_39,
	b_ram_data_in_bus_23,
	b_ram_data_in_bus_7,
	b_ram_data_in_bus_55,
	b_ram_data_in_bus_38,
	b_ram_data_in_bus_22,
	b_ram_data_in_bus_6,
	b_ram_data_in_bus_54,
	b_ram_data_in_bus_35,
	b_ram_data_in_bus_19,
	b_ram_data_in_bus_3,
	b_ram_data_in_bus_51,
	b_ram_data_in_bus_36,
	b_ram_data_in_bus_20,
	b_ram_data_in_bus_4,
	b_ram_data_in_bus_52,
	b_ram_data_in_bus_37,
	b_ram_data_in_bus_21,
	b_ram_data_in_bus_5,
	b_ram_data_in_bus_53,
	b_ram_data_in_bus_34,
	b_ram_data_in_bus_18,
	b_ram_data_in_bus_2,
	b_ram_data_in_bus_50,
	b_ram_data_in_bus_24,
	b_ram_data_in_bus_8,
	b_ram_data_in_bus_56,
	b_ram_data_in_bus_40,
	b_ram_data_in_bus_25,
	b_ram_data_in_bus_9,
	b_ram_data_in_bus_57,
	b_ram_data_in_bus_41,
	b_ram_data_in_bus_0,
	b_ram_data_in_bus_48,
	b_ram_data_in_bus_32,
	b_ram_data_in_bus_16,
	b_ram_data_in_bus_1,
	b_ram_data_in_bus_49,
	b_ram_data_in_bus_33,
	b_ram_data_in_bus_17,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_141;
output 	q_b_142;
output 	q_b_143;
output 	q_b_13;
output 	q_b_131;
output 	q_b_132;
output 	q_b_133;
output 	q_b_10;
output 	q_b_101;
output 	q_b_102;
output 	q_b_103;
output 	q_b_11;
output 	q_b_111;
output 	q_b_112;
output 	q_b_113;
output 	q_b_12;
output 	q_b_121;
output 	q_b_122;
output 	q_b_123;
output 	q_b_15;
output 	q_b_151;
output 	q_b_152;
output 	q_b_153;
output 	q_b_7;
output 	q_b_71;
output 	q_b_72;
output 	q_b_73;
output 	q_b_6;
output 	q_b_61;
output 	q_b_62;
output 	q_b_63;
output 	q_b_3;
output 	q_b_31;
output 	q_b_32;
output 	q_b_33;
output 	q_b_4;
output 	q_b_41;
output 	q_b_42;
output 	q_b_43;
output 	q_b_5;
output 	q_b_51;
output 	q_b_52;
output 	q_b_53;
output 	q_b_2;
output 	q_b_21;
output 	q_b_22;
output 	q_b_23;
output 	q_b_8;
output 	q_b_81;
output 	q_b_82;
output 	q_b_83;
output 	q_b_9;
output 	q_b_91;
output 	q_b_92;
output 	q_b_93;
output 	q_b_0;
output 	q_b_01;
output 	q_b_02;
output 	q_b_03;
output 	q_b_1;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
input 	wren_b_1;
input 	b_ram_data_in_bus_46;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_9;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_9;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wren_b_2;
input 	b_ram_data_in_bus_30;
input 	wraddress_b_bus_12;
input 	wraddress_b_bus_5;
input 	rdaddress_b_bus_12;
input 	rdaddress_b_bus_5;
input 	wren_b_3;
input 	b_ram_data_in_bus_14;
input 	wraddress_b_bus_1;
input 	rdaddress_b_bus_1;
input 	wren_b_0;
input 	b_ram_data_in_bus_62;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_45;
input 	b_ram_data_in_bus_29;
input 	b_ram_data_in_bus_13;
input 	b_ram_data_in_bus_61;
input 	b_ram_data_in_bus_42;
input 	b_ram_data_in_bus_26;
input 	b_ram_data_in_bus_10;
input 	b_ram_data_in_bus_58;
input 	b_ram_data_in_bus_43;
input 	b_ram_data_in_bus_27;
input 	b_ram_data_in_bus_11;
input 	b_ram_data_in_bus_59;
input 	b_ram_data_in_bus_44;
input 	b_ram_data_in_bus_28;
input 	b_ram_data_in_bus_12;
input 	b_ram_data_in_bus_60;
input 	b_ram_data_in_bus_47;
input 	b_ram_data_in_bus_31;
input 	b_ram_data_in_bus_15;
input 	b_ram_data_in_bus_63;
input 	b_ram_data_in_bus_39;
input 	b_ram_data_in_bus_23;
input 	b_ram_data_in_bus_7;
input 	b_ram_data_in_bus_55;
input 	b_ram_data_in_bus_38;
input 	b_ram_data_in_bus_22;
input 	b_ram_data_in_bus_6;
input 	b_ram_data_in_bus_54;
input 	b_ram_data_in_bus_35;
input 	b_ram_data_in_bus_19;
input 	b_ram_data_in_bus_3;
input 	b_ram_data_in_bus_51;
input 	b_ram_data_in_bus_36;
input 	b_ram_data_in_bus_20;
input 	b_ram_data_in_bus_4;
input 	b_ram_data_in_bus_52;
input 	b_ram_data_in_bus_37;
input 	b_ram_data_in_bus_21;
input 	b_ram_data_in_bus_5;
input 	b_ram_data_in_bus_53;
input 	b_ram_data_in_bus_34;
input 	b_ram_data_in_bus_18;
input 	b_ram_data_in_bus_2;
input 	b_ram_data_in_bus_50;
input 	b_ram_data_in_bus_24;
input 	b_ram_data_in_bus_8;
input 	b_ram_data_in_bus_56;
input 	b_ram_data_in_bus_40;
input 	b_ram_data_in_bus_25;
input 	b_ram_data_in_bus_9;
input 	b_ram_data_in_bus_57;
input 	b_ram_data_in_bus_41;
input 	b_ram_data_in_bus_0;
input 	b_ram_data_in_bus_48;
input 	b_ram_data_in_bus_32;
input 	b_ram_data_in_bus_16;
input 	b_ram_data_in_bus_1;
input 	b_ram_data_in_bus_49;
input 	b_ram_data_in_bus_33;
input 	b_ram_data_in_bus_17;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_asj_fft_data_ram_12 \gen_rams:0:dat_A (
	.q_b_14(q_b_143),
	.q_b_13(q_b_133),
	.q_b_10(q_b_103),
	.q_b_11(q_b_113),
	.q_b_12(q_b_123),
	.q_b_15(q_b_153),
	.q_b_7(q_b_73),
	.q_b_6(q_b_63),
	.q_b_3(q_b_33),
	.q_b_4(q_b_43),
	.q_b_5(q_b_53),
	.q_b_2(q_b_23),
	.q_b_8(q_b_82),
	.q_b_9(q_b_92),
	.q_b_0(q_b_01),
	.q_b_1(q_b_16),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.wraddress_b_bus_12(wraddress_b_bus_12),
	.rdaddress_b_bus_12(rdaddress_b_bus_12),
	.wren_b_0(wren_b_0),
	.b_ram_data_in_bus_62(b_ram_data_in_bus_62),
	.wraddress_b_bus_13(wraddress_b_bus_13),
	.rdaddress_b_bus_13(rdaddress_b_bus_13),
	.b_ram_data_in_bus_61(b_ram_data_in_bus_61),
	.b_ram_data_in_bus_58(b_ram_data_in_bus_58),
	.b_ram_data_in_bus_59(b_ram_data_in_bus_59),
	.b_ram_data_in_bus_60(b_ram_data_in_bus_60),
	.b_ram_data_in_bus_63(b_ram_data_in_bus_63),
	.b_ram_data_in_bus_55(b_ram_data_in_bus_55),
	.b_ram_data_in_bus_54(b_ram_data_in_bus_54),
	.b_ram_data_in_bus_51(b_ram_data_in_bus_51),
	.b_ram_data_in_bus_52(b_ram_data_in_bus_52),
	.b_ram_data_in_bus_53(b_ram_data_in_bus_53),
	.b_ram_data_in_bus_50(b_ram_data_in_bus_50),
	.b_ram_data_in_bus_56(b_ram_data_in_bus_56),
	.b_ram_data_in_bus_57(b_ram_data_in_bus_57),
	.b_ram_data_in_bus_48(b_ram_data_in_bus_48),
	.b_ram_data_in_bus_49(b_ram_data_in_bus_49),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

IFFT_asj_fft_data_ram_13 \gen_rams:1:dat_A (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_83),
	.q_b_9(q_b_93),
	.q_b_0(q_b_02),
	.q_b_1(q_b_17),
	.wren_b_1(wren_b_1),
	.b_ram_data_in_bus_46(b_ram_data_in_bus_46),
	.wraddress_b_bus_0(wraddress_b_bus_0),
	.wraddress_b_bus_9(wraddress_b_bus_9),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_0(rdaddress_b_bus_0),
	.rdaddress_b_bus_9(rdaddress_b_bus_9),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.b_ram_data_in_bus_45(b_ram_data_in_bus_45),
	.b_ram_data_in_bus_42(b_ram_data_in_bus_42),
	.b_ram_data_in_bus_43(b_ram_data_in_bus_43),
	.b_ram_data_in_bus_44(b_ram_data_in_bus_44),
	.b_ram_data_in_bus_47(b_ram_data_in_bus_47),
	.b_ram_data_in_bus_39(b_ram_data_in_bus_39),
	.b_ram_data_in_bus_38(b_ram_data_in_bus_38),
	.b_ram_data_in_bus_35(b_ram_data_in_bus_35),
	.b_ram_data_in_bus_36(b_ram_data_in_bus_36),
	.b_ram_data_in_bus_37(b_ram_data_in_bus_37),
	.b_ram_data_in_bus_34(b_ram_data_in_bus_34),
	.b_ram_data_in_bus_40(b_ram_data_in_bus_40),
	.b_ram_data_in_bus_41(b_ram_data_in_bus_41),
	.b_ram_data_in_bus_32(b_ram_data_in_bus_32),
	.b_ram_data_in_bus_33(b_ram_data_in_bus_33),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

IFFT_asj_fft_data_ram_15 \gen_rams:3:dat_A (
	.q_b_14(q_b_142),
	.q_b_13(q_b_132),
	.q_b_10(q_b_102),
	.q_b_11(q_b_112),
	.q_b_12(q_b_122),
	.q_b_15(q_b_152),
	.q_b_7(q_b_72),
	.q_b_6(q_b_62),
	.q_b_3(q_b_32),
	.q_b_4(q_b_42),
	.q_b_5(q_b_52),
	.q_b_2(q_b_22),
	.q_b_8(q_b_81),
	.q_b_9(q_b_91),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_b_bus_0(wraddress_b_bus_0),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_0(rdaddress_b_bus_0),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.wren_b_3(wren_b_3),
	.b_ram_data_in_bus_14(b_ram_data_in_bus_14),
	.wraddress_b_bus_1(wraddress_b_bus_1),
	.rdaddress_b_bus_1(rdaddress_b_bus_1),
	.b_ram_data_in_bus_13(b_ram_data_in_bus_13),
	.b_ram_data_in_bus_10(b_ram_data_in_bus_10),
	.b_ram_data_in_bus_11(b_ram_data_in_bus_11),
	.b_ram_data_in_bus_12(b_ram_data_in_bus_12),
	.b_ram_data_in_bus_15(b_ram_data_in_bus_15),
	.b_ram_data_in_bus_7(b_ram_data_in_bus_7),
	.b_ram_data_in_bus_6(b_ram_data_in_bus_6),
	.b_ram_data_in_bus_3(b_ram_data_in_bus_3),
	.b_ram_data_in_bus_4(b_ram_data_in_bus_4),
	.b_ram_data_in_bus_5(b_ram_data_in_bus_5),
	.b_ram_data_in_bus_2(b_ram_data_in_bus_2),
	.b_ram_data_in_bus_8(b_ram_data_in_bus_8),
	.b_ram_data_in_bus_9(b_ram_data_in_bus_9),
	.b_ram_data_in_bus_0(b_ram_data_in_bus_0),
	.b_ram_data_in_bus_1(b_ram_data_in_bus_1),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

IFFT_asj_fft_data_ram_14 \gen_rams:2:dat_A (
	.q_b_14(q_b_141),
	.q_b_13(q_b_131),
	.q_b_10(q_b_101),
	.q_b_11(q_b_111),
	.q_b_12(q_b_121),
	.q_b_15(q_b_151),
	.q_b_7(q_b_71),
	.q_b_6(q_b_61),
	.q_b_3(q_b_31),
	.q_b_4(q_b_41),
	.q_b_5(q_b_51),
	.q_b_2(q_b_21),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_03),
	.q_b_1(q_b_18),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.wren_b_2(wren_b_2),
	.b_ram_data_in_bus_30(b_ram_data_in_bus_30),
	.wraddress_b_bus_12(wraddress_b_bus_12),
	.wraddress_b_bus_5(wraddress_b_bus_5),
	.rdaddress_b_bus_12(rdaddress_b_bus_12),
	.rdaddress_b_bus_5(rdaddress_b_bus_5),
	.b_ram_data_in_bus_29(b_ram_data_in_bus_29),
	.b_ram_data_in_bus_26(b_ram_data_in_bus_26),
	.b_ram_data_in_bus_27(b_ram_data_in_bus_27),
	.b_ram_data_in_bus_28(b_ram_data_in_bus_28),
	.b_ram_data_in_bus_31(b_ram_data_in_bus_31),
	.b_ram_data_in_bus_23(b_ram_data_in_bus_23),
	.b_ram_data_in_bus_22(b_ram_data_in_bus_22),
	.b_ram_data_in_bus_19(b_ram_data_in_bus_19),
	.b_ram_data_in_bus_20(b_ram_data_in_bus_20),
	.b_ram_data_in_bus_21(b_ram_data_in_bus_21),
	.b_ram_data_in_bus_18(b_ram_data_in_bus_18),
	.b_ram_data_in_bus_24(b_ram_data_in_bus_24),
	.b_ram_data_in_bus_25(b_ram_data_in_bus_25),
	.b_ram_data_in_bus_16(b_ram_data_in_bus_16),
	.b_ram_data_in_bus_17(b_ram_data_in_bus_17),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_asj_fft_data_ram_12 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wraddress_b_bus_12,
	rdaddress_b_bus_12,
	wren_b_0,
	b_ram_data_in_bus_62,
	wraddress_b_bus_13,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_61,
	b_ram_data_in_bus_58,
	b_ram_data_in_bus_59,
	b_ram_data_in_bus_60,
	b_ram_data_in_bus_63,
	b_ram_data_in_bus_55,
	b_ram_data_in_bus_54,
	b_ram_data_in_bus_51,
	b_ram_data_in_bus_52,
	b_ram_data_in_bus_53,
	b_ram_data_in_bus_50,
	b_ram_data_in_bus_56,
	b_ram_data_in_bus_57,
	b_ram_data_in_bus_48,
	b_ram_data_in_bus_49,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wraddress_b_bus_12;
input 	rdaddress_b_bus_12;
input 	wren_b_0;
input 	b_ram_data_in_bus_62;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_61;
input 	b_ram_data_in_bus_58;
input 	b_ram_data_in_bus_59;
input 	b_ram_data_in_bus_60;
input 	b_ram_data_in_bus_63;
input 	b_ram_data_in_bus_55;
input 	b_ram_data_in_bus_54;
input 	b_ram_data_in_bus_51;
input 	b_ram_data_in_bus_52;
input 	b_ram_data_in_bus_53;
input 	b_ram_data_in_bus_50;
input 	b_ram_data_in_bus_56;
input 	b_ram_data_in_bus_57;
input 	b_ram_data_in_bus_48;
input 	b_ram_data_in_bus_49;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_12 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.wraddress_b_bus_12(wraddress_b_bus_12),
	.rdaddress_b_bus_12(rdaddress_b_bus_12),
	.wren_b_0(wren_b_0),
	.b_ram_data_in_bus_62(b_ram_data_in_bus_62),
	.wraddress_b_bus_13(wraddress_b_bus_13),
	.rdaddress_b_bus_13(rdaddress_b_bus_13),
	.b_ram_data_in_bus_61(b_ram_data_in_bus_61),
	.b_ram_data_in_bus_58(b_ram_data_in_bus_58),
	.b_ram_data_in_bus_59(b_ram_data_in_bus_59),
	.b_ram_data_in_bus_60(b_ram_data_in_bus_60),
	.b_ram_data_in_bus_63(b_ram_data_in_bus_63),
	.b_ram_data_in_bus_55(b_ram_data_in_bus_55),
	.b_ram_data_in_bus_54(b_ram_data_in_bus_54),
	.b_ram_data_in_bus_51(b_ram_data_in_bus_51),
	.b_ram_data_in_bus_52(b_ram_data_in_bus_52),
	.b_ram_data_in_bus_53(b_ram_data_in_bus_53),
	.b_ram_data_in_bus_50(b_ram_data_in_bus_50),
	.b_ram_data_in_bus_56(b_ram_data_in_bus_56),
	.b_ram_data_in_bus_57(b_ram_data_in_bus_57),
	.b_ram_data_in_bus_48(b_ram_data_in_bus_48),
	.b_ram_data_in_bus_49(b_ram_data_in_bus_49),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_12 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wraddress_b_bus_12,
	rdaddress_b_bus_12,
	wren_b_0,
	b_ram_data_in_bus_62,
	wraddress_b_bus_13,
	rdaddress_b_bus_13,
	b_ram_data_in_bus_61,
	b_ram_data_in_bus_58,
	b_ram_data_in_bus_59,
	b_ram_data_in_bus_60,
	b_ram_data_in_bus_63,
	b_ram_data_in_bus_55,
	b_ram_data_in_bus_54,
	b_ram_data_in_bus_51,
	b_ram_data_in_bus_52,
	b_ram_data_in_bus_53,
	b_ram_data_in_bus_50,
	b_ram_data_in_bus_56,
	b_ram_data_in_bus_57,
	b_ram_data_in_bus_48,
	b_ram_data_in_bus_49,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wraddress_b_bus_12;
input 	rdaddress_b_bus_12;
input 	wren_b_0;
input 	b_ram_data_in_bus_62;
input 	wraddress_b_bus_13;
input 	rdaddress_b_bus_13;
input 	b_ram_data_in_bus_61;
input 	b_ram_data_in_bus_58;
input 	b_ram_data_in_bus_59;
input 	b_ram_data_in_bus_60;
input 	b_ram_data_in_bus_63;
input 	b_ram_data_in_bus_55;
input 	b_ram_data_in_bus_54;
input 	b_ram_data_in_bus_51;
input 	b_ram_data_in_bus_52;
input 	b_ram_data_in_bus_53;
input 	b_ram_data_in_bus_50;
input 	b_ram_data_in_bus_56;
input 	b_ram_data_in_bus_57;
input 	b_ram_data_in_bus_48;
input 	b_ram_data_in_bus_49;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_19 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({wraddress_b_bus_11,wraddress_b_bus_10,wraddress_b_bus_13,wraddress_b_bus_12}),
	.address_b({rdaddress_b_bus_11,rdaddress_b_bus_10,rdaddress_b_bus_13,rdaddress_b_bus_12}),
	.wren_a(wren_b_0),
	.data_a({b_ram_data_in_bus_63,b_ram_data_in_bus_62,b_ram_data_in_bus_61,b_ram_data_in_bus_60,b_ram_data_in_bus_59,b_ram_data_in_bus_58,b_ram_data_in_bus_57,b_ram_data_in_bus_56,b_ram_data_in_bus_55,b_ram_data_in_bus_54,b_ram_data_in_bus_53,b_ram_data_in_bus_52,
b_ram_data_in_bus_51,b_ram_data_in_bus_50,b_ram_data_in_bus_49,b_ram_data_in_bus_48}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_19 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_12 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_12 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:0:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_13 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wren_b_1,
	b_ram_data_in_bus_46,
	wraddress_b_bus_0,
	wraddress_b_bus_9,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_0,
	rdaddress_b_bus_9,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	b_ram_data_in_bus_45,
	b_ram_data_in_bus_42,
	b_ram_data_in_bus_43,
	b_ram_data_in_bus_44,
	b_ram_data_in_bus_47,
	b_ram_data_in_bus_39,
	b_ram_data_in_bus_38,
	b_ram_data_in_bus_35,
	b_ram_data_in_bus_36,
	b_ram_data_in_bus_37,
	b_ram_data_in_bus_34,
	b_ram_data_in_bus_40,
	b_ram_data_in_bus_41,
	b_ram_data_in_bus_32,
	b_ram_data_in_bus_33,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wren_b_1;
input 	b_ram_data_in_bus_46;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_9;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_9;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	b_ram_data_in_bus_45;
input 	b_ram_data_in_bus_42;
input 	b_ram_data_in_bus_43;
input 	b_ram_data_in_bus_44;
input 	b_ram_data_in_bus_47;
input 	b_ram_data_in_bus_39;
input 	b_ram_data_in_bus_38;
input 	b_ram_data_in_bus_35;
input 	b_ram_data_in_bus_36;
input 	b_ram_data_in_bus_37;
input 	b_ram_data_in_bus_34;
input 	b_ram_data_in_bus_40;
input 	b_ram_data_in_bus_41;
input 	b_ram_data_in_bus_32;
input 	b_ram_data_in_bus_33;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_13 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wren_b_1(wren_b_1),
	.b_ram_data_in_bus_46(b_ram_data_in_bus_46),
	.wraddress_b_bus_0(wraddress_b_bus_0),
	.wraddress_b_bus_9(wraddress_b_bus_9),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_0(rdaddress_b_bus_0),
	.rdaddress_b_bus_9(rdaddress_b_bus_9),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.b_ram_data_in_bus_45(b_ram_data_in_bus_45),
	.b_ram_data_in_bus_42(b_ram_data_in_bus_42),
	.b_ram_data_in_bus_43(b_ram_data_in_bus_43),
	.b_ram_data_in_bus_44(b_ram_data_in_bus_44),
	.b_ram_data_in_bus_47(b_ram_data_in_bus_47),
	.b_ram_data_in_bus_39(b_ram_data_in_bus_39),
	.b_ram_data_in_bus_38(b_ram_data_in_bus_38),
	.b_ram_data_in_bus_35(b_ram_data_in_bus_35),
	.b_ram_data_in_bus_36(b_ram_data_in_bus_36),
	.b_ram_data_in_bus_37(b_ram_data_in_bus_37),
	.b_ram_data_in_bus_34(b_ram_data_in_bus_34),
	.b_ram_data_in_bus_40(b_ram_data_in_bus_40),
	.b_ram_data_in_bus_41(b_ram_data_in_bus_41),
	.b_ram_data_in_bus_32(b_ram_data_in_bus_32),
	.b_ram_data_in_bus_33(b_ram_data_in_bus_33),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_13 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wren_b_1,
	b_ram_data_in_bus_46,
	wraddress_b_bus_0,
	wraddress_b_bus_9,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_0,
	rdaddress_b_bus_9,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	b_ram_data_in_bus_45,
	b_ram_data_in_bus_42,
	b_ram_data_in_bus_43,
	b_ram_data_in_bus_44,
	b_ram_data_in_bus_47,
	b_ram_data_in_bus_39,
	b_ram_data_in_bus_38,
	b_ram_data_in_bus_35,
	b_ram_data_in_bus_36,
	b_ram_data_in_bus_37,
	b_ram_data_in_bus_34,
	b_ram_data_in_bus_40,
	b_ram_data_in_bus_41,
	b_ram_data_in_bus_32,
	b_ram_data_in_bus_33,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wren_b_1;
input 	b_ram_data_in_bus_46;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_9;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_9;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	b_ram_data_in_bus_45;
input 	b_ram_data_in_bus_42;
input 	b_ram_data_in_bus_43;
input 	b_ram_data_in_bus_44;
input 	b_ram_data_in_bus_47;
input 	b_ram_data_in_bus_39;
input 	b_ram_data_in_bus_38;
input 	b_ram_data_in_bus_35;
input 	b_ram_data_in_bus_36;
input 	b_ram_data_in_bus_37;
input 	b_ram_data_in_bus_34;
input 	b_ram_data_in_bus_40;
input 	b_ram_data_in_bus_41;
input 	b_ram_data_in_bus_32;
input 	b_ram_data_in_bus_33;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_20 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(wren_b_1),
	.data_a({b_ram_data_in_bus_47,b_ram_data_in_bus_46,b_ram_data_in_bus_45,b_ram_data_in_bus_44,b_ram_data_in_bus_43,b_ram_data_in_bus_42,b_ram_data_in_bus_41,b_ram_data_in_bus_40,b_ram_data_in_bus_39,b_ram_data_in_bus_38,b_ram_data_in_bus_37,b_ram_data_in_bus_36,
b_ram_data_in_bus_35,b_ram_data_in_bus_34,b_ram_data_in_bus_33,b_ram_data_in_bus_32}),
	.address_a({wraddress_b_bus_11,wraddress_b_bus_10,wraddress_b_bus_9,wraddress_b_bus_0}),
	.address_b({rdaddress_b_bus_11,rdaddress_b_bus_10,rdaddress_b_bus_9,rdaddress_b_bus_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_20 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[15:0] data_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_13 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_13 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[15:0] data_a;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:1:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_14 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wren_b_2,
	b_ram_data_in_bus_30,
	wraddress_b_bus_12,
	wraddress_b_bus_5,
	rdaddress_b_bus_12,
	rdaddress_b_bus_5,
	b_ram_data_in_bus_29,
	b_ram_data_in_bus_26,
	b_ram_data_in_bus_27,
	b_ram_data_in_bus_28,
	b_ram_data_in_bus_31,
	b_ram_data_in_bus_23,
	b_ram_data_in_bus_22,
	b_ram_data_in_bus_19,
	b_ram_data_in_bus_20,
	b_ram_data_in_bus_21,
	b_ram_data_in_bus_18,
	b_ram_data_in_bus_24,
	b_ram_data_in_bus_25,
	b_ram_data_in_bus_16,
	b_ram_data_in_bus_17,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wren_b_2;
input 	b_ram_data_in_bus_30;
input 	wraddress_b_bus_12;
input 	wraddress_b_bus_5;
input 	rdaddress_b_bus_12;
input 	rdaddress_b_bus_5;
input 	b_ram_data_in_bus_29;
input 	b_ram_data_in_bus_26;
input 	b_ram_data_in_bus_27;
input 	b_ram_data_in_bus_28;
input 	b_ram_data_in_bus_31;
input 	b_ram_data_in_bus_23;
input 	b_ram_data_in_bus_22;
input 	b_ram_data_in_bus_19;
input 	b_ram_data_in_bus_20;
input 	b_ram_data_in_bus_21;
input 	b_ram_data_in_bus_18;
input 	b_ram_data_in_bus_24;
input 	b_ram_data_in_bus_25;
input 	b_ram_data_in_bus_16;
input 	b_ram_data_in_bus_17;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_14 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.wren_b_2(wren_b_2),
	.b_ram_data_in_bus_30(b_ram_data_in_bus_30),
	.wraddress_b_bus_12(wraddress_b_bus_12),
	.wraddress_b_bus_5(wraddress_b_bus_5),
	.rdaddress_b_bus_12(rdaddress_b_bus_12),
	.rdaddress_b_bus_5(rdaddress_b_bus_5),
	.b_ram_data_in_bus_29(b_ram_data_in_bus_29),
	.b_ram_data_in_bus_26(b_ram_data_in_bus_26),
	.b_ram_data_in_bus_27(b_ram_data_in_bus_27),
	.b_ram_data_in_bus_28(b_ram_data_in_bus_28),
	.b_ram_data_in_bus_31(b_ram_data_in_bus_31),
	.b_ram_data_in_bus_23(b_ram_data_in_bus_23),
	.b_ram_data_in_bus_22(b_ram_data_in_bus_22),
	.b_ram_data_in_bus_19(b_ram_data_in_bus_19),
	.b_ram_data_in_bus_20(b_ram_data_in_bus_20),
	.b_ram_data_in_bus_21(b_ram_data_in_bus_21),
	.b_ram_data_in_bus_18(b_ram_data_in_bus_18),
	.b_ram_data_in_bus_24(b_ram_data_in_bus_24),
	.b_ram_data_in_bus_25(b_ram_data_in_bus_25),
	.b_ram_data_in_bus_16(b_ram_data_in_bus_16),
	.b_ram_data_in_bus_17(b_ram_data_in_bus_17),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_14 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wren_b_2,
	b_ram_data_in_bus_30,
	wraddress_b_bus_12,
	wraddress_b_bus_5,
	rdaddress_b_bus_12,
	rdaddress_b_bus_5,
	b_ram_data_in_bus_29,
	b_ram_data_in_bus_26,
	b_ram_data_in_bus_27,
	b_ram_data_in_bus_28,
	b_ram_data_in_bus_31,
	b_ram_data_in_bus_23,
	b_ram_data_in_bus_22,
	b_ram_data_in_bus_19,
	b_ram_data_in_bus_20,
	b_ram_data_in_bus_21,
	b_ram_data_in_bus_18,
	b_ram_data_in_bus_24,
	b_ram_data_in_bus_25,
	b_ram_data_in_bus_16,
	b_ram_data_in_bus_17,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wren_b_2;
input 	b_ram_data_in_bus_30;
input 	wraddress_b_bus_12;
input 	wraddress_b_bus_5;
input 	rdaddress_b_bus_12;
input 	rdaddress_b_bus_5;
input 	b_ram_data_in_bus_29;
input 	b_ram_data_in_bus_26;
input 	b_ram_data_in_bus_27;
input 	b_ram_data_in_bus_28;
input 	b_ram_data_in_bus_31;
input 	b_ram_data_in_bus_23;
input 	b_ram_data_in_bus_22;
input 	b_ram_data_in_bus_19;
input 	b_ram_data_in_bus_20;
input 	b_ram_data_in_bus_21;
input 	b_ram_data_in_bus_18;
input 	b_ram_data_in_bus_24;
input 	b_ram_data_in_bus_25;
input 	b_ram_data_in_bus_16;
input 	b_ram_data_in_bus_17;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_21 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({wraddress_b_bus_11,wraddress_b_bus_10,wraddress_b_bus_5,wraddress_b_bus_12}),
	.address_b({rdaddress_b_bus_11,rdaddress_b_bus_10,rdaddress_b_bus_5,rdaddress_b_bus_12}),
	.wren_a(wren_b_2),
	.data_a({b_ram_data_in_bus_31,b_ram_data_in_bus_30,b_ram_data_in_bus_29,b_ram_data_in_bus_28,b_ram_data_in_bus_27,b_ram_data_in_bus_26,b_ram_data_in_bus_25,b_ram_data_in_bus_24,b_ram_data_in_bus_23,b_ram_data_in_bus_22,b_ram_data_in_bus_21,b_ram_data_in_bus_20,
b_ram_data_in_bus_19,b_ram_data_in_bus_18,b_ram_data_in_bus_17,b_ram_data_in_bus_16}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_21 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_14 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_14 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:2:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_data_ram_15 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_b_bus_0,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_0,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wren_b_3,
	b_ram_data_in_bus_14,
	wraddress_b_bus_1,
	rdaddress_b_bus_1,
	b_ram_data_in_bus_13,
	b_ram_data_in_bus_10,
	b_ram_data_in_bus_11,
	b_ram_data_in_bus_12,
	b_ram_data_in_bus_15,
	b_ram_data_in_bus_7,
	b_ram_data_in_bus_6,
	b_ram_data_in_bus_3,
	b_ram_data_in_bus_4,
	b_ram_data_in_bus_5,
	b_ram_data_in_bus_2,
	b_ram_data_in_bus_8,
	b_ram_data_in_bus_9,
	b_ram_data_in_bus_0,
	b_ram_data_in_bus_1,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wren_b_3;
input 	b_ram_data_in_bus_14;
input 	wraddress_b_bus_1;
input 	rdaddress_b_bus_1;
input 	b_ram_data_in_bus_13;
input 	b_ram_data_in_bus_10;
input 	b_ram_data_in_bus_11;
input 	b_ram_data_in_bus_12;
input 	b_ram_data_in_bus_15;
input 	b_ram_data_in_bus_7;
input 	b_ram_data_in_bus_6;
input 	b_ram_data_in_bus_3;
input 	b_ram_data_in_bus_4;
input 	b_ram_data_in_bus_5;
input 	b_ram_data_in_bus_2;
input 	b_ram_data_in_bus_8;
input 	b_ram_data_in_bus_9;
input 	b_ram_data_in_bus_0;
input 	b_ram_data_in_bus_1;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altera_fft_dual_port_ram_15 \gen_M4K:ram_component (
	.q_b_14(q_b_14),
	.q_b_13(q_b_13),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_15(q_b_15),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_2(q_b_2),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.wraddress_b_bus_0(wraddress_b_bus_0),
	.wraddress_b_bus_10(wraddress_b_bus_10),
	.wraddress_b_bus_11(wraddress_b_bus_11),
	.rdaddress_b_bus_0(rdaddress_b_bus_0),
	.rdaddress_b_bus_10(rdaddress_b_bus_10),
	.rdaddress_b_bus_11(rdaddress_b_bus_11),
	.wren_b_3(wren_b_3),
	.b_ram_data_in_bus_14(b_ram_data_in_bus_14),
	.wraddress_b_bus_1(wraddress_b_bus_1),
	.rdaddress_b_bus_1(rdaddress_b_bus_1),
	.b_ram_data_in_bus_13(b_ram_data_in_bus_13),
	.b_ram_data_in_bus_10(b_ram_data_in_bus_10),
	.b_ram_data_in_bus_11(b_ram_data_in_bus_11),
	.b_ram_data_in_bus_12(b_ram_data_in_bus_12),
	.b_ram_data_in_bus_15(b_ram_data_in_bus_15),
	.b_ram_data_in_bus_7(b_ram_data_in_bus_7),
	.b_ram_data_in_bus_6(b_ram_data_in_bus_6),
	.b_ram_data_in_bus_3(b_ram_data_in_bus_3),
	.b_ram_data_in_bus_4(b_ram_data_in_bus_4),
	.b_ram_data_in_bus_5(b_ram_data_in_bus_5),
	.b_ram_data_in_bus_2(b_ram_data_in_bus_2),
	.b_ram_data_in_bus_8(b_ram_data_in_bus_8),
	.b_ram_data_in_bus_9(b_ram_data_in_bus_9),
	.b_ram_data_in_bus_0(b_ram_data_in_bus_0),
	.b_ram_data_in_bus_1(b_ram_data_in_bus_1),
	.global_clock_enable(global_clock_enable),
	.clk(clk));

endmodule

module IFFT_altera_fft_dual_port_ram_15 (
	q_b_14,
	q_b_13,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_15,
	q_b_7,
	q_b_6,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_2,
	q_b_8,
	q_b_9,
	q_b_0,
	q_b_1,
	wraddress_b_bus_0,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_0,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	wren_b_3,
	b_ram_data_in_bus_14,
	wraddress_b_bus_1,
	rdaddress_b_bus_1,
	b_ram_data_in_bus_13,
	b_ram_data_in_bus_10,
	b_ram_data_in_bus_11,
	b_ram_data_in_bus_12,
	b_ram_data_in_bus_15,
	b_ram_data_in_bus_7,
	b_ram_data_in_bus_6,
	b_ram_data_in_bus_3,
	b_ram_data_in_bus_4,
	b_ram_data_in_bus_5,
	b_ram_data_in_bus_2,
	b_ram_data_in_bus_8,
	b_ram_data_in_bus_9,
	b_ram_data_in_bus_0,
	b_ram_data_in_bus_1,
	global_clock_enable,
	clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_14;
output 	q_b_13;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_15;
output 	q_b_7;
output 	q_b_6;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_2;
output 	q_b_8;
output 	q_b_9;
output 	q_b_0;
output 	q_b_1;
input 	wraddress_b_bus_0;
input 	wraddress_b_bus_10;
input 	wraddress_b_bus_11;
input 	rdaddress_b_bus_0;
input 	rdaddress_b_bus_10;
input 	rdaddress_b_bus_11;
input 	wren_b_3;
input 	b_ram_data_in_bus_14;
input 	wraddress_b_bus_1;
input 	rdaddress_b_bus_1;
input 	b_ram_data_in_bus_13;
input 	b_ram_data_in_bus_10;
input 	b_ram_data_in_bus_11;
input 	b_ram_data_in_bus_12;
input 	b_ram_data_in_bus_15;
input 	b_ram_data_in_bus_7;
input 	b_ram_data_in_bus_6;
input 	b_ram_data_in_bus_3;
input 	b_ram_data_in_bus_4;
input 	b_ram_data_in_bus_5;
input 	b_ram_data_in_bus_2;
input 	b_ram_data_in_bus_8;
input 	b_ram_data_in_bus_9;
input 	b_ram_data_in_bus_0;
input 	b_ram_data_in_bus_1;
input 	global_clock_enable;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_22 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({wraddress_b_bus_11,wraddress_b_bus_10,wraddress_b_bus_1,wraddress_b_bus_0}),
	.address_b({rdaddress_b_bus_11,rdaddress_b_bus_10,rdaddress_b_bus_1,rdaddress_b_bus_0}),
	.wren_a(wren_b_3),
	.data_a({b_ram_data_in_bus_15,b_ram_data_in_bus_14,b_ram_data_in_bus_13,b_ram_data_in_bus_12,b_ram_data_in_bus_11,b_ram_data_in_bus_10,b_ram_data_in_bus_9,b_ram_data_in_bus_8,b_ram_data_in_bus_7,b_ram_data_in_bus_6,b_ram_data_in_bus_5,b_ram_data_in_bus_4,b_ram_data_in_bus_3,
b_ram_data_in_bus_2,b_ram_data_in_bus_1,b_ram_data_in_bus_0}),
	.clocken0(global_clock_enable),
	.clock0(clk));

endmodule

module IFFT_altsyncram_22 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_altsyncram_j304_15 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clocken0(clocken0),
	.clock0(clock0));

endmodule

module IFFT_altsyncram_j304_15 (
	q_b,
	address_a,
	address_b,
	wren_a,
	data_a,
	clocken0,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[3:0] address_a;
input 	[3:0] address_b;
input 	wren_a;
input 	[15:0] data_a;
input 	clocken0;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_4dp_ram:dat_B|asj_fft_data_ram:\\gen_rams:3:dat_A|altera_fft_dual_port_ram:\\gen_M4K:ram_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_j304:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_asj_fft_bfp_ctrl (
	tdl_arr_4,
	tdl_arr_11,
	global_clock_enable,
	blk_exp_0,
	blk_exp_1,
	blk_exp_2,
	blk_exp_3,
	blk_exp_4,
	blk_exp_5,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	lut_out_tmp_0,
	lut_out_tmp_1,
	lut_out_tmp_2,
	en_slb,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	tdl_arr_4;
input 	tdl_arr_11;
input 	global_clock_enable;
output 	blk_exp_0;
output 	blk_exp_1;
output 	blk_exp_2;
output 	blk_exp_3;
output 	blk_exp_4;
output 	blk_exp_5;
output 	slb_last_0;
output 	slb_last_1;
output 	slb_last_2;
input 	lut_out_tmp_0;
input 	lut_out_tmp_1;
input 	lut_out_tmp_2;
input 	en_slb;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass2|tdl_arr[0]~q ;
wire \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ;
wire \Add0~1_sumout ;
wire \blk_exp_acc[0]~0_combout ;
wire \blk_exp_acc[0]~1_combout ;
wire \blk_exp_acc[0]~q ;
wire \blk_exp~0_combout ;
wire \blk_exp[0]~1_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \blk_exp_acc[1]~q ;
wire \blk_exp~2_combout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \blk_exp_acc[2]~q ;
wire \blk_exp~3_combout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \blk_exp_acc[3]~q ;
wire \blk_exp~4_combout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \blk_exp_acc[4]~q ;
wire \blk_exp~5_combout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \blk_exp_acc[5]~q ;
wire \blk_exp~6_combout ;
wire \slb_last~0_combout ;
wire \slb_last[2]~1_combout ;
wire \slb_last~2_combout ;
wire \slb_last~3_combout ;


IFFT_asj_fft_tdl_bit_rst_1 \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass2 (
	.tdl_arr_0(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass2|tdl_arr[0]~q ),
	.tdl_arr_8(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_tdl_bit_rst \gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass (
	.tdl_arr_8(\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ),
	.global_clock_enable(global_clock_enable),
	.en_slb(en_slb),
	.clk(clk),
	.reset_n(reset_n));

dffeas \blk_exp[0] (
	.clk(clk),
	.d(\blk_exp~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_0),
	.prn(vcc));
defparam \blk_exp[0] .is_wysiwyg = "true";
defparam \blk_exp[0] .power_up = "low";

dffeas \blk_exp[1] (
	.clk(clk),
	.d(\blk_exp~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_1),
	.prn(vcc));
defparam \blk_exp[1] .is_wysiwyg = "true";
defparam \blk_exp[1] .power_up = "low";

dffeas \blk_exp[2] (
	.clk(clk),
	.d(\blk_exp~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_2),
	.prn(vcc));
defparam \blk_exp[2] .is_wysiwyg = "true";
defparam \blk_exp[2] .power_up = "low";

dffeas \blk_exp[3] (
	.clk(clk),
	.d(\blk_exp~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_3),
	.prn(vcc));
defparam \blk_exp[3] .is_wysiwyg = "true";
defparam \blk_exp[3] .power_up = "low";

dffeas \blk_exp[4] (
	.clk(clk),
	.d(\blk_exp~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_4),
	.prn(vcc));
defparam \blk_exp[4] .is_wysiwyg = "true";
defparam \blk_exp[4] .power_up = "low";

dffeas \blk_exp[5] (
	.clk(clk),
	.d(\blk_exp~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\blk_exp[0]~1_combout ),
	.q(blk_exp_5),
	.prn(vcc));
defparam \blk_exp[5] .is_wysiwyg = "true";
defparam \blk_exp[5] .power_up = "low";

dffeas \slb_last[0] (
	.clk(clk),
	.d(\slb_last~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~1_combout ),
	.q(slb_last_0),
	.prn(vcc));
defparam \slb_last[0] .is_wysiwyg = "true";
defparam \slb_last[0] .power_up = "low";

dffeas \slb_last[1] (
	.clk(clk),
	.d(\slb_last~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~1_combout ),
	.q(slb_last_1),
	.prn(vcc));
defparam \slb_last[1] .is_wysiwyg = "true";
defparam \slb_last[1] .power_up = "low";

dffeas \slb_last[2] (
	.clk(clk),
	.d(\slb_last~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\slb_last[2]~1_combout ),
	.q(slb_last_2),
	.prn(vcc));
defparam \slb_last[2] .is_wysiwyg = "true";
defparam \slb_last[2] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\blk_exp_acc[0]~q ),
	.datae(gnd),
	.dataf(!slb_last_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \blk_exp_acc[0]~0 (
	.dataa(!reset_n),
	.datab(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass2|tdl_arr[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp_acc[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp_acc[0]~0 .extended_lut = "off";
defparam \blk_exp_acc[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \blk_exp_acc[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \blk_exp_acc[0]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass2|tdl_arr[0]~q ),
	.datad(!tdl_arr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp_acc[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp_acc[0]~1 .extended_lut = "off";
defparam \blk_exp_acc[0]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \blk_exp_acc[0]~1 .shared_arith = "off";

dffeas \blk_exp_acc[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~0_combout ),
	.ena(\blk_exp_acc[0]~1_combout ),
	.q(\blk_exp_acc[0]~q ),
	.prn(vcc));
defparam \blk_exp_acc[0] .is_wysiwyg = "true";
defparam \blk_exp_acc[0] .power_up = "low";

cyclonev_lcell_comb \blk_exp~0 (
	.dataa(!reset_n),
	.datab(!\blk_exp_acc[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp~0 .extended_lut = "off";
defparam \blk_exp~0 .lut_mask = 64'h7777777777777777;
defparam \blk_exp~0 .shared_arith = "off";

cyclonev_lcell_comb \blk_exp[0]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass2|tdl_arr[0]~q ),
	.datad(!tdl_arr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp[0]~1 .extended_lut = "off";
defparam \blk_exp[0]~1 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \blk_exp[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\blk_exp_acc[1]~q ),
	.datae(gnd),
	.dataf(!slb_last_1),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \blk_exp_acc[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~0_combout ),
	.ena(\blk_exp_acc[0]~1_combout ),
	.q(\blk_exp_acc[1]~q ),
	.prn(vcc));
defparam \blk_exp_acc[1] .is_wysiwyg = "true";
defparam \blk_exp_acc[1] .power_up = "low";

cyclonev_lcell_comb \blk_exp~2 (
	.dataa(!reset_n),
	.datab(!\blk_exp_acc[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp~2 .extended_lut = "off";
defparam \blk_exp~2 .lut_mask = 64'h7777777777777777;
defparam \blk_exp~2 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\blk_exp_acc[2]~q ),
	.datae(gnd),
	.dataf(!slb_last_2),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \blk_exp_acc[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~0_combout ),
	.ena(\blk_exp_acc[0]~1_combout ),
	.q(\blk_exp_acc[2]~q ),
	.prn(vcc));
defparam \blk_exp_acc[2] .is_wysiwyg = "true";
defparam \blk_exp_acc[2] .power_up = "low";

cyclonev_lcell_comb \blk_exp~3 (
	.dataa(!reset_n),
	.datab(!\blk_exp_acc[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp~3 .extended_lut = "off";
defparam \blk_exp~3 .lut_mask = 64'h7777777777777777;
defparam \blk_exp~3 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\blk_exp_acc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \blk_exp_acc[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~0_combout ),
	.ena(\blk_exp_acc[0]~1_combout ),
	.q(\blk_exp_acc[3]~q ),
	.prn(vcc));
defparam \blk_exp_acc[3] .is_wysiwyg = "true";
defparam \blk_exp_acc[3] .power_up = "low";

cyclonev_lcell_comb \blk_exp~4 (
	.dataa(!reset_n),
	.datab(!\blk_exp_acc[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp~4 .extended_lut = "off";
defparam \blk_exp~4 .lut_mask = 64'h7777777777777777;
defparam \blk_exp~4 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\blk_exp_acc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \blk_exp_acc[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~0_combout ),
	.ena(\blk_exp_acc[0]~1_combout ),
	.q(\blk_exp_acc[4]~q ),
	.prn(vcc));
defparam \blk_exp_acc[4] .is_wysiwyg = "true";
defparam \blk_exp_acc[4] .power_up = "low";

cyclonev_lcell_comb \blk_exp~5 (
	.dataa(!reset_n),
	.datab(!\blk_exp_acc[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp~5 .extended_lut = "off";
defparam \blk_exp~5 .lut_mask = 64'h7777777777777777;
defparam \blk_exp~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\blk_exp_acc[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \blk_exp_acc[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\blk_exp_acc[0]~0_combout ),
	.ena(\blk_exp_acc[0]~1_combout ),
	.q(\blk_exp_acc[5]~q ),
	.prn(vcc));
defparam \blk_exp_acc[5] .is_wysiwyg = "true";
defparam \blk_exp_acc[5] .power_up = "low";

cyclonev_lcell_comb \blk_exp~6 (
	.dataa(!reset_n),
	.datab(!\blk_exp_acc[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_exp~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_exp~6 .extended_lut = "off";
defparam \blk_exp~6 .lut_mask = 64'h7777777777777777;
defparam \blk_exp~6 .shared_arith = "off";

cyclonev_lcell_comb \slb_last~0 (
	.dataa(!reset_n),
	.datab(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ),
	.datac(!lut_out_tmp_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_last~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_last~0 .extended_lut = "off";
defparam \slb_last~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \slb_last~0 .shared_arith = "off";

cyclonev_lcell_comb \slb_last[2]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ),
	.datad(!tdl_arr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_last[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_last[2]~1 .extended_lut = "off";
defparam \slb_last[2]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \slb_last[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \slb_last~2 (
	.dataa(!reset_n),
	.datab(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ),
	.datac(!lut_out_tmp_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_last~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_last~2 .extended_lut = "off";
defparam \slb_last~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \slb_last~2 .shared_arith = "off";

cyclonev_lcell_comb \slb_last~3 (
	.dataa(!reset_n),
	.datab(!\gen_quad_str_ctrl:gen_se_bfp:gen_4bit_accum:gen_disc:delay_next_pass|tdl_arr[8]~q ),
	.datac(!lut_out_tmp_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_last~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_last~3 .extended_lut = "off";
defparam \slb_last~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \slb_last~3 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl_bit_rst (
	tdl_arr_8,
	global_clock_enable,
	en_slb,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_8;
input 	global_clock_enable;
input 	en_slb;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;


dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_8),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(en_slb),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_bit_rst_1 (
	tdl_arr_0,
	tdl_arr_8,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_0;
input 	tdl_arr_8;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(tdl_arr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module IFFT_asj_fft_cnt_ctrl (
	ram_block6a0,
	ram_block6a1,
	data_rdy_vec_10,
	q_b_14,
	q_b_141,
	q_b_142,
	q_b_143,
	q_b_144,
	q_b_145,
	q_b_146,
	q_b_147,
	q_b_13,
	q_b_131,
	q_b_132,
	q_b_133,
	q_b_134,
	q_b_135,
	q_b_136,
	q_b_137,
	q_b_10,
	q_b_101,
	q_b_102,
	q_b_103,
	q_b_104,
	q_b_105,
	q_b_106,
	q_b_107,
	q_b_11,
	q_b_111,
	q_b_112,
	q_b_113,
	q_b_114,
	q_b_115,
	q_b_116,
	q_b_117,
	q_b_12,
	q_b_121,
	q_b_122,
	q_b_123,
	q_b_124,
	q_b_125,
	q_b_126,
	q_b_127,
	q_b_15,
	q_b_151,
	q_b_152,
	q_b_153,
	q_b_154,
	q_b_155,
	q_b_156,
	q_b_157,
	q_b_7,
	q_b_71,
	q_b_72,
	q_b_73,
	q_b_74,
	q_b_75,
	q_b_76,
	q_b_77,
	q_b_6,
	q_b_61,
	q_b_62,
	q_b_63,
	q_b_64,
	q_b_65,
	q_b_66,
	q_b_67,
	q_b_3,
	q_b_31,
	q_b_32,
	q_b_33,
	q_b_34,
	q_b_35,
	q_b_36,
	q_b_37,
	q_b_4,
	q_b_41,
	q_b_42,
	q_b_43,
	q_b_44,
	q_b_45,
	q_b_46,
	q_b_47,
	q_b_5,
	q_b_51,
	q_b_52,
	q_b_53,
	q_b_54,
	q_b_55,
	q_b_56,
	q_b_57,
	q_b_2,
	q_b_21,
	q_b_22,
	q_b_23,
	q_b_24,
	q_b_25,
	q_b_26,
	q_b_27,
	q_b_8,
	q_b_81,
	q_b_82,
	q_b_83,
	q_b_84,
	q_b_85,
	q_b_86,
	q_b_87,
	q_b_9,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_94,
	q_b_95,
	q_b_96,
	q_b_97,
	q_b_0,
	q_b_01,
	q_b_02,
	q_b_03,
	q_b_04,
	q_b_05,
	q_b_06,
	q_b_07,
	q_b_1,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_110,
	q_b_118,
	q_b_119,
	b_ram_data_in_bus_46,
	wraddress_b_bus_0,
	wraddress_b_bus_9,
	wraddress_b_bus_10,
	wraddress_b_bus_11,
	rdaddress_b_bus_0,
	rdaddress_b_bus_9,
	rdaddress_b_bus_10,
	rdaddress_b_bus_11,
	a_ram_data_in_bus_46,
	wraddress_a_bus_0,
	wraddress_a_bus_9,
	wraddress_a_bus_10,
	wraddress_a_bus_11,
	rdaddress_a_bus_0,
	rdaddress_a_bus_9,
	rdaddress_a_bus_10,
	rdaddress_a_bus_11,
	b_ram_data_in_bus_30,
	wraddress_b_bus_12,
	wraddress_b_bus_5,
	rdaddress_b_bus_12,
	rdaddress_b_bus_5,
	a_ram_data_in_bus_30,
	wraddress_a_bus_12,
	wraddress_a_bus_5,
	rdaddress_a_bus_12,
	rdaddress_a_bus_5,
	b_ram_data_in_bus_14,
	wraddress_b_bus_1,
	rdaddress_b_bus_1,
	a_ram_data_in_bus_14,
	wraddress_a_bus_1,
	rdaddress_a_bus_1,
	b_ram_data_in_bus_62,
	wraddress_b_bus_13,
	rdaddress_b_bus_13,
	a_ram_data_in_bus_62,
	wraddress_a_bus_13,
	rdaddress_a_bus_13,
	b_ram_data_in_bus_45,
	a_ram_data_in_bus_45,
	b_ram_data_in_bus_29,
	a_ram_data_in_bus_29,
	b_ram_data_in_bus_13,
	a_ram_data_in_bus_13,
	b_ram_data_in_bus_61,
	a_ram_data_in_bus_61,
	b_ram_data_in_bus_42,
	a_ram_data_in_bus_42,
	b_ram_data_in_bus_26,
	a_ram_data_in_bus_26,
	b_ram_data_in_bus_10,
	a_ram_data_in_bus_10,
	b_ram_data_in_bus_58,
	a_ram_data_in_bus_58,
	b_ram_data_in_bus_43,
	a_ram_data_in_bus_43,
	b_ram_data_in_bus_27,
	a_ram_data_in_bus_27,
	b_ram_data_in_bus_11,
	a_ram_data_in_bus_11,
	b_ram_data_in_bus_59,
	a_ram_data_in_bus_59,
	b_ram_data_in_bus_44,
	a_ram_data_in_bus_44,
	b_ram_data_in_bus_28,
	a_ram_data_in_bus_28,
	b_ram_data_in_bus_12,
	a_ram_data_in_bus_12,
	b_ram_data_in_bus_60,
	a_ram_data_in_bus_60,
	b_ram_data_in_bus_47,
	a_ram_data_in_bus_47,
	b_ram_data_in_bus_31,
	a_ram_data_in_bus_31,
	b_ram_data_in_bus_15,
	a_ram_data_in_bus_15,
	b_ram_data_in_bus_63,
	a_ram_data_in_bus_63,
	b_ram_data_in_bus_39,
	a_ram_data_in_bus_39,
	b_ram_data_in_bus_23,
	a_ram_data_in_bus_23,
	b_ram_data_in_bus_7,
	a_ram_data_in_bus_7,
	b_ram_data_in_bus_55,
	a_ram_data_in_bus_55,
	b_ram_data_in_bus_38,
	a_ram_data_in_bus_38,
	b_ram_data_in_bus_22,
	a_ram_data_in_bus_22,
	b_ram_data_in_bus_6,
	a_ram_data_in_bus_6,
	b_ram_data_in_bus_54,
	a_ram_data_in_bus_54,
	b_ram_data_in_bus_35,
	a_ram_data_in_bus_35,
	b_ram_data_in_bus_19,
	a_ram_data_in_bus_19,
	b_ram_data_in_bus_3,
	a_ram_data_in_bus_3,
	b_ram_data_in_bus_51,
	a_ram_data_in_bus_51,
	b_ram_data_in_bus_36,
	a_ram_data_in_bus_36,
	b_ram_data_in_bus_20,
	a_ram_data_in_bus_20,
	b_ram_data_in_bus_4,
	a_ram_data_in_bus_4,
	b_ram_data_in_bus_52,
	a_ram_data_in_bus_52,
	b_ram_data_in_bus_37,
	a_ram_data_in_bus_37,
	b_ram_data_in_bus_21,
	a_ram_data_in_bus_21,
	b_ram_data_in_bus_5,
	a_ram_data_in_bus_5,
	b_ram_data_in_bus_53,
	a_ram_data_in_bus_53,
	b_ram_data_in_bus_34,
	a_ram_data_in_bus_34,
	b_ram_data_in_bus_18,
	a_ram_data_in_bus_18,
	b_ram_data_in_bus_2,
	a_ram_data_in_bus_2,
	b_ram_data_in_bus_50,
	a_ram_data_in_bus_50,
	b_ram_data_in_bus_24,
	a_ram_data_in_bus_24,
	b_ram_data_in_bus_8,
	a_ram_data_in_bus_8,
	b_ram_data_in_bus_56,
	a_ram_data_in_bus_56,
	b_ram_data_in_bus_40,
	a_ram_data_in_bus_40,
	b_ram_data_in_bus_25,
	a_ram_data_in_bus_25,
	b_ram_data_in_bus_9,
	a_ram_data_in_bus_9,
	b_ram_data_in_bus_57,
	a_ram_data_in_bus_57,
	b_ram_data_in_bus_41,
	a_ram_data_in_bus_41,
	b_ram_data_in_bus_0,
	a_ram_data_in_bus_0,
	b_ram_data_in_bus_48,
	a_ram_data_in_bus_48,
	b_ram_data_in_bus_32,
	a_ram_data_in_bus_32,
	b_ram_data_in_bus_16,
	a_ram_data_in_bus_16,
	b_ram_data_in_bus_1,
	a_ram_data_in_bus_1,
	b_ram_data_in_bus_49,
	a_ram_data_in_bus_49,
	b_ram_data_in_bus_33,
	a_ram_data_in_bus_33,
	b_ram_data_in_bus_17,
	a_ram_data_in_bus_17,
	data_in_r_6,
	wr_address_i_int_0,
	wr_address_i_int_1,
	wr_address_i_int_2,
	wr_address_i_int_3,
	data_in_r_5,
	data_in_r_2,
	data_in_r_3,
	data_in_r_4,
	data_in_r_7,
	data_in_i_7,
	data_in_i_6,
	data_in_i_3,
	data_in_i_4,
	data_in_i_5,
	data_in_i_2,
	data_in_r_0,
	data_in_r_1,
	data_in_i_0,
	data_in_i_1,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_2_0,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_1,
	ram_in_reg_1_1,
	ram_in_reg_2_2,
	ram_in_reg_1_2,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_5,
	ram_in_reg_2_6,
	ram_in_reg_3_3,
	ram_in_reg_3_0,
	ram_in_reg_3_1,
	ram_in_reg_3_2,
	ram_in_reg_3_7,
	ram_in_reg_3_4,
	ram_in_reg_3_5,
	ram_in_reg_3_6,
	ram_in_reg_4_3,
	ram_in_reg_4_0,
	ram_in_reg_4_1,
	ram_in_reg_4_2,
	ram_in_reg_4_7,
	ram_in_reg_4_4,
	ram_in_reg_4_5,
	ram_in_reg_4_6,
	ram_in_reg_5_3,
	ram_in_reg_5_0,
	ram_in_reg_5_1,
	ram_in_reg_5_2,
	ram_in_reg_5_7,
	ram_in_reg_5_4,
	ram_in_reg_5_5,
	ram_in_reg_5_6,
	ram_in_reg_6_3,
	ram_in_reg_6_0,
	ram_in_reg_6_1,
	ram_in_reg_6_2,
	ram_in_reg_6_7,
	ram_in_reg_6_4,
	ram_in_reg_6_5,
	ram_in_reg_6_6,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_1,
	ram_in_reg_7_2,
	ram_in_reg_7_7,
	ram_in_reg_7_4,
	ram_in_reg_7_5,
	ram_in_reg_7_6,
	ram_in_reg_2_01,
	ram_in_reg_3_01,
	ram_in_reg_1_31,
	ram_in_reg_1_01,
	ram_in_reg_1_11,
	ram_in_reg_1_21,
	ram_in_reg_1_7,
	ram_in_reg_1_4,
	ram_in_reg_1_5,
	ram_in_reg_1_6,
	ram_in_reg_0_01,
	ram_in_reg_0_11,
	ram_in_reg_1_32,
	ram_in_reg_1_12,
	ram_in_reg_1_22,
	ram_in_reg_1_02,
	ram_in_reg_0_3,
	ram_in_reg_0_02,
	ram_in_reg_0_12,
	ram_in_reg_0_2,
	ram_in_reg_0_7,
	ram_in_reg_0_4,
	ram_in_reg_0_5,
	ram_in_reg_0_6,
	ram_data_out1_14,
	ram_data_out2_14,
	ram_data_out3_14,
	ram_data_out0_14,
	ram_data_out1_13,
	ram_data_out2_13,
	ram_data_out3_13,
	ram_data_out0_13,
	ram_data_out1_10,
	ram_data_out2_10,
	ram_data_out3_10,
	ram_data_out0_10,
	ram_data_out1_11,
	ram_data_out2_11,
	ram_data_out3_11,
	ram_data_out0_11,
	ram_data_out1_12,
	ram_data_out2_12,
	ram_data_out3_12,
	ram_data_out0_12,
	ram_data_out1_15,
	ram_data_out2_15,
	ram_data_out3_15,
	ram_data_out0_15,
	ram_data_out1_7,
	ram_data_out2_7,
	ram_data_out3_7,
	ram_data_out0_7,
	ram_data_out1_6,
	ram_data_out2_6,
	ram_data_out3_6,
	ram_data_out0_6,
	ram_data_out1_3,
	ram_data_out2_3,
	ram_data_out3_3,
	ram_data_out0_3,
	ram_data_out1_4,
	ram_data_out2_4,
	ram_data_out3_4,
	ram_data_out0_4,
	ram_data_out1_5,
	ram_data_out2_5,
	ram_data_out3_5,
	ram_data_out0_5,
	ram_data_out1_2,
	ram_data_out2_2,
	ram_data_out3_2,
	ram_data_out0_2,
	ram_data_out2_8,
	ram_data_out3_8,
	ram_data_out0_8,
	ram_data_out1_8,
	ram_data_out2_9,
	ram_data_out3_9,
	ram_data_out0_9,
	ram_data_out1_9,
	ram_data_out3_0,
	ram_data_out0_0,
	ram_data_out1_0,
	ram_data_out2_0,
	ram_data_out3_1,
	ram_data_out0_1,
	ram_data_out1_1,
	ram_data_out2_1,
	ram_a_not_b_vec_10,
	ram_a_not_b_vec_1,
	sel_anb_addr,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ram_block6a0;
input 	ram_block6a1;
input 	data_rdy_vec_10;
input 	q_b_14;
input 	q_b_141;
input 	q_b_142;
input 	q_b_143;
input 	q_b_144;
input 	q_b_145;
input 	q_b_146;
input 	q_b_147;
input 	q_b_13;
input 	q_b_131;
input 	q_b_132;
input 	q_b_133;
input 	q_b_134;
input 	q_b_135;
input 	q_b_136;
input 	q_b_137;
input 	q_b_10;
input 	q_b_101;
input 	q_b_102;
input 	q_b_103;
input 	q_b_104;
input 	q_b_105;
input 	q_b_106;
input 	q_b_107;
input 	q_b_11;
input 	q_b_111;
input 	q_b_112;
input 	q_b_113;
input 	q_b_114;
input 	q_b_115;
input 	q_b_116;
input 	q_b_117;
input 	q_b_12;
input 	q_b_121;
input 	q_b_122;
input 	q_b_123;
input 	q_b_124;
input 	q_b_125;
input 	q_b_126;
input 	q_b_127;
input 	q_b_15;
input 	q_b_151;
input 	q_b_152;
input 	q_b_153;
input 	q_b_154;
input 	q_b_155;
input 	q_b_156;
input 	q_b_157;
input 	q_b_7;
input 	q_b_71;
input 	q_b_72;
input 	q_b_73;
input 	q_b_74;
input 	q_b_75;
input 	q_b_76;
input 	q_b_77;
input 	q_b_6;
input 	q_b_61;
input 	q_b_62;
input 	q_b_63;
input 	q_b_64;
input 	q_b_65;
input 	q_b_66;
input 	q_b_67;
input 	q_b_3;
input 	q_b_31;
input 	q_b_32;
input 	q_b_33;
input 	q_b_34;
input 	q_b_35;
input 	q_b_36;
input 	q_b_37;
input 	q_b_4;
input 	q_b_41;
input 	q_b_42;
input 	q_b_43;
input 	q_b_44;
input 	q_b_45;
input 	q_b_46;
input 	q_b_47;
input 	q_b_5;
input 	q_b_51;
input 	q_b_52;
input 	q_b_53;
input 	q_b_54;
input 	q_b_55;
input 	q_b_56;
input 	q_b_57;
input 	q_b_2;
input 	q_b_21;
input 	q_b_22;
input 	q_b_23;
input 	q_b_24;
input 	q_b_25;
input 	q_b_26;
input 	q_b_27;
input 	q_b_8;
input 	q_b_81;
input 	q_b_82;
input 	q_b_83;
input 	q_b_84;
input 	q_b_85;
input 	q_b_86;
input 	q_b_87;
input 	q_b_9;
input 	q_b_91;
input 	q_b_92;
input 	q_b_93;
input 	q_b_94;
input 	q_b_95;
input 	q_b_96;
input 	q_b_97;
input 	q_b_0;
input 	q_b_01;
input 	q_b_02;
input 	q_b_03;
input 	q_b_04;
input 	q_b_05;
input 	q_b_06;
input 	q_b_07;
input 	q_b_1;
input 	q_b_16;
input 	q_b_17;
input 	q_b_18;
input 	q_b_19;
input 	q_b_110;
input 	q_b_118;
input 	q_b_119;
output 	b_ram_data_in_bus_46;
output 	wraddress_b_bus_0;
output 	wraddress_b_bus_9;
output 	wraddress_b_bus_10;
output 	wraddress_b_bus_11;
output 	rdaddress_b_bus_0;
output 	rdaddress_b_bus_9;
output 	rdaddress_b_bus_10;
output 	rdaddress_b_bus_11;
output 	a_ram_data_in_bus_46;
output 	wraddress_a_bus_0;
output 	wraddress_a_bus_9;
output 	wraddress_a_bus_10;
output 	wraddress_a_bus_11;
output 	rdaddress_a_bus_0;
output 	rdaddress_a_bus_9;
output 	rdaddress_a_bus_10;
output 	rdaddress_a_bus_11;
output 	b_ram_data_in_bus_30;
output 	wraddress_b_bus_12;
output 	wraddress_b_bus_5;
output 	rdaddress_b_bus_12;
output 	rdaddress_b_bus_5;
output 	a_ram_data_in_bus_30;
output 	wraddress_a_bus_12;
output 	wraddress_a_bus_5;
output 	rdaddress_a_bus_12;
output 	rdaddress_a_bus_5;
output 	b_ram_data_in_bus_14;
output 	wraddress_b_bus_1;
output 	rdaddress_b_bus_1;
output 	a_ram_data_in_bus_14;
output 	wraddress_a_bus_1;
output 	rdaddress_a_bus_1;
output 	b_ram_data_in_bus_62;
output 	wraddress_b_bus_13;
output 	rdaddress_b_bus_13;
output 	a_ram_data_in_bus_62;
output 	wraddress_a_bus_13;
output 	rdaddress_a_bus_13;
output 	b_ram_data_in_bus_45;
output 	a_ram_data_in_bus_45;
output 	b_ram_data_in_bus_29;
output 	a_ram_data_in_bus_29;
output 	b_ram_data_in_bus_13;
output 	a_ram_data_in_bus_13;
output 	b_ram_data_in_bus_61;
output 	a_ram_data_in_bus_61;
output 	b_ram_data_in_bus_42;
output 	a_ram_data_in_bus_42;
output 	b_ram_data_in_bus_26;
output 	a_ram_data_in_bus_26;
output 	b_ram_data_in_bus_10;
output 	a_ram_data_in_bus_10;
output 	b_ram_data_in_bus_58;
output 	a_ram_data_in_bus_58;
output 	b_ram_data_in_bus_43;
output 	a_ram_data_in_bus_43;
output 	b_ram_data_in_bus_27;
output 	a_ram_data_in_bus_27;
output 	b_ram_data_in_bus_11;
output 	a_ram_data_in_bus_11;
output 	b_ram_data_in_bus_59;
output 	a_ram_data_in_bus_59;
output 	b_ram_data_in_bus_44;
output 	a_ram_data_in_bus_44;
output 	b_ram_data_in_bus_28;
output 	a_ram_data_in_bus_28;
output 	b_ram_data_in_bus_12;
output 	a_ram_data_in_bus_12;
output 	b_ram_data_in_bus_60;
output 	a_ram_data_in_bus_60;
output 	b_ram_data_in_bus_47;
output 	a_ram_data_in_bus_47;
output 	b_ram_data_in_bus_31;
output 	a_ram_data_in_bus_31;
output 	b_ram_data_in_bus_15;
output 	a_ram_data_in_bus_15;
output 	b_ram_data_in_bus_63;
output 	a_ram_data_in_bus_63;
output 	b_ram_data_in_bus_39;
output 	a_ram_data_in_bus_39;
output 	b_ram_data_in_bus_23;
output 	a_ram_data_in_bus_23;
output 	b_ram_data_in_bus_7;
output 	a_ram_data_in_bus_7;
output 	b_ram_data_in_bus_55;
output 	a_ram_data_in_bus_55;
output 	b_ram_data_in_bus_38;
output 	a_ram_data_in_bus_38;
output 	b_ram_data_in_bus_22;
output 	a_ram_data_in_bus_22;
output 	b_ram_data_in_bus_6;
output 	a_ram_data_in_bus_6;
output 	b_ram_data_in_bus_54;
output 	a_ram_data_in_bus_54;
output 	b_ram_data_in_bus_35;
output 	a_ram_data_in_bus_35;
output 	b_ram_data_in_bus_19;
output 	a_ram_data_in_bus_19;
output 	b_ram_data_in_bus_3;
output 	a_ram_data_in_bus_3;
output 	b_ram_data_in_bus_51;
output 	a_ram_data_in_bus_51;
output 	b_ram_data_in_bus_36;
output 	a_ram_data_in_bus_36;
output 	b_ram_data_in_bus_20;
output 	a_ram_data_in_bus_20;
output 	b_ram_data_in_bus_4;
output 	a_ram_data_in_bus_4;
output 	b_ram_data_in_bus_52;
output 	a_ram_data_in_bus_52;
output 	b_ram_data_in_bus_37;
output 	a_ram_data_in_bus_37;
output 	b_ram_data_in_bus_21;
output 	a_ram_data_in_bus_21;
output 	b_ram_data_in_bus_5;
output 	a_ram_data_in_bus_5;
output 	b_ram_data_in_bus_53;
output 	a_ram_data_in_bus_53;
output 	b_ram_data_in_bus_34;
output 	a_ram_data_in_bus_34;
output 	b_ram_data_in_bus_18;
output 	a_ram_data_in_bus_18;
output 	b_ram_data_in_bus_2;
output 	a_ram_data_in_bus_2;
output 	b_ram_data_in_bus_50;
output 	a_ram_data_in_bus_50;
output 	b_ram_data_in_bus_24;
output 	a_ram_data_in_bus_24;
output 	b_ram_data_in_bus_8;
output 	a_ram_data_in_bus_8;
output 	b_ram_data_in_bus_56;
output 	a_ram_data_in_bus_56;
output 	b_ram_data_in_bus_40;
output 	a_ram_data_in_bus_40;
output 	b_ram_data_in_bus_25;
output 	a_ram_data_in_bus_25;
output 	b_ram_data_in_bus_9;
output 	a_ram_data_in_bus_9;
output 	b_ram_data_in_bus_57;
output 	a_ram_data_in_bus_57;
output 	b_ram_data_in_bus_41;
output 	a_ram_data_in_bus_41;
output 	b_ram_data_in_bus_0;
output 	a_ram_data_in_bus_0;
output 	b_ram_data_in_bus_48;
output 	a_ram_data_in_bus_48;
output 	b_ram_data_in_bus_32;
output 	a_ram_data_in_bus_32;
output 	b_ram_data_in_bus_16;
output 	a_ram_data_in_bus_16;
output 	b_ram_data_in_bus_1;
output 	a_ram_data_in_bus_1;
output 	b_ram_data_in_bus_49;
output 	a_ram_data_in_bus_49;
output 	b_ram_data_in_bus_33;
output 	a_ram_data_in_bus_33;
output 	b_ram_data_in_bus_17;
output 	a_ram_data_in_bus_17;
input 	data_in_r_6;
input 	wr_address_i_int_0;
input 	wr_address_i_int_1;
input 	wr_address_i_int_2;
input 	wr_address_i_int_3;
input 	data_in_r_5;
input 	data_in_r_2;
input 	data_in_r_3;
input 	data_in_r_4;
input 	data_in_r_7;
input 	data_in_i_7;
input 	data_in_i_6;
input 	data_in_i_3;
input 	data_in_i_4;
input 	data_in_i_5;
input 	data_in_i_2;
input 	data_in_r_0;
input 	data_in_r_1;
input 	data_in_i_0;
input 	data_in_i_1;
input 	global_clock_enable;
input 	ram_in_reg_2_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_3;
input 	ram_in_reg_2_0;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_2_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_2_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_6;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_0;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_2;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_4;
input 	ram_in_reg_3_5;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_0;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_2;
input 	ram_in_reg_4_7;
input 	ram_in_reg_4_4;
input 	ram_in_reg_4_5;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_0;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_2;
input 	ram_in_reg_5_7;
input 	ram_in_reg_5_4;
input 	ram_in_reg_5_5;
input 	ram_in_reg_5_6;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_0;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_2;
input 	ram_in_reg_6_7;
input 	ram_in_reg_6_4;
input 	ram_in_reg_6_5;
input 	ram_in_reg_6_6;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_7;
input 	ram_in_reg_7_4;
input 	ram_in_reg_7_5;
input 	ram_in_reg_7_6;
input 	ram_in_reg_2_01;
input 	ram_in_reg_3_01;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_01;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_4;
input 	ram_in_reg_1_5;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_32;
input 	ram_in_reg_1_12;
input 	ram_in_reg_1_22;
input 	ram_in_reg_1_02;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_02;
input 	ram_in_reg_0_12;
input 	ram_in_reg_0_2;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_4;
input 	ram_in_reg_0_5;
input 	ram_in_reg_0_6;
output 	ram_data_out1_14;
output 	ram_data_out2_14;
output 	ram_data_out3_14;
output 	ram_data_out0_14;
output 	ram_data_out1_13;
output 	ram_data_out2_13;
output 	ram_data_out3_13;
output 	ram_data_out0_13;
output 	ram_data_out1_10;
output 	ram_data_out2_10;
output 	ram_data_out3_10;
output 	ram_data_out0_10;
output 	ram_data_out1_11;
output 	ram_data_out2_11;
output 	ram_data_out3_11;
output 	ram_data_out0_11;
output 	ram_data_out1_12;
output 	ram_data_out2_12;
output 	ram_data_out3_12;
output 	ram_data_out0_12;
output 	ram_data_out1_15;
output 	ram_data_out2_15;
output 	ram_data_out3_15;
output 	ram_data_out0_15;
output 	ram_data_out1_7;
output 	ram_data_out2_7;
output 	ram_data_out3_7;
output 	ram_data_out0_7;
output 	ram_data_out1_6;
output 	ram_data_out2_6;
output 	ram_data_out3_6;
output 	ram_data_out0_6;
output 	ram_data_out1_3;
output 	ram_data_out2_3;
output 	ram_data_out3_3;
output 	ram_data_out0_3;
output 	ram_data_out1_4;
output 	ram_data_out2_4;
output 	ram_data_out3_4;
output 	ram_data_out0_4;
output 	ram_data_out1_5;
output 	ram_data_out2_5;
output 	ram_data_out3_5;
output 	ram_data_out0_5;
output 	ram_data_out1_2;
output 	ram_data_out2_2;
output 	ram_data_out3_2;
output 	ram_data_out0_2;
output 	ram_data_out2_8;
output 	ram_data_out3_8;
output 	ram_data_out0_8;
output 	ram_data_out1_8;
output 	ram_data_out2_9;
output 	ram_data_out3_9;
output 	ram_data_out0_9;
output 	ram_data_out1_9;
output 	ram_data_out3_0;
output 	ram_data_out0_0;
output 	ram_data_out1_0;
output 	ram_data_out2_0;
output 	ram_data_out3_1;
output 	ram_data_out0_1;
output 	ram_data_out1_1;
output 	ram_data_out2_1;
input 	ram_a_not_b_vec_10;
input 	ram_a_not_b_vec_1;
input 	sel_anb_addr;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_data_out1~0_combout ;
wire \ram_data_out2~0_combout ;
wire \ram_data_out3~0_combout ;
wire \ram_data_out0~0_combout ;
wire \ram_data_out1~1_combout ;
wire \ram_data_out2~1_combout ;
wire \ram_data_out3~1_combout ;
wire \ram_data_out0~1_combout ;
wire \ram_data_out1~2_combout ;
wire \ram_data_out2~2_combout ;
wire \ram_data_out3~2_combout ;
wire \ram_data_out0~2_combout ;
wire \ram_data_out1~3_combout ;
wire \ram_data_out2~3_combout ;
wire \ram_data_out3~3_combout ;
wire \ram_data_out0~3_combout ;
wire \ram_data_out1~4_combout ;
wire \ram_data_out2~4_combout ;
wire \ram_data_out3~4_combout ;
wire \ram_data_out0~4_combout ;
wire \ram_data_out1~5_combout ;
wire \ram_data_out2~5_combout ;
wire \ram_data_out3~5_combout ;
wire \ram_data_out0~5_combout ;
wire \ram_data_out1~6_combout ;
wire \ram_data_out2~6_combout ;
wire \ram_data_out3~6_combout ;
wire \ram_data_out0~6_combout ;
wire \ram_data_out1~7_combout ;
wire \ram_data_out2~7_combout ;
wire \ram_data_out3~7_combout ;
wire \ram_data_out0~7_combout ;
wire \ram_data_out1~8_combout ;
wire \ram_data_out2~8_combout ;
wire \ram_data_out3~8_combout ;
wire \ram_data_out0~8_combout ;
wire \ram_data_out1~9_combout ;
wire \ram_data_out2~9_combout ;
wire \ram_data_out3~9_combout ;
wire \ram_data_out0~9_combout ;
wire \ram_data_out1~10_combout ;
wire \ram_data_out2~10_combout ;
wire \ram_data_out3~10_combout ;
wire \ram_data_out0~10_combout ;
wire \ram_data_out1~11_combout ;
wire \ram_data_out2~11_combout ;
wire \ram_data_out3~11_combout ;
wire \ram_data_out0~11_combout ;
wire \ram_data_out2~12_combout ;
wire \ram_data_out3~12_combout ;
wire \ram_data_out0~12_combout ;
wire \ram_data_out1~12_combout ;
wire \ram_data_out2~13_combout ;
wire \ram_data_out3~13_combout ;
wire \ram_data_out0~13_combout ;
wire \ram_data_out1~13_combout ;
wire \ram_data_out3~14_combout ;
wire \ram_data_out0~14_combout ;
wire \ram_data_out1~14_combout ;
wire \ram_data_out2~14_combout ;
wire \ram_data_out3~15_combout ;
wire \ram_data_out0~15_combout ;
wire \ram_data_out1~15_combout ;
wire \ram_data_out2~15_combout ;


dffeas \b_ram_data_in_bus[46] (
	.clk(clk),
	.d(ram_in_reg_6_1),
	.asdata(data_in_r_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_46),
	.prn(vcc));
defparam \b_ram_data_in_bus[46] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[46] .power_up = "low";

dffeas \wraddress_b_bus[0] (
	.clk(clk),
	.d(ram_in_reg_0_1),
	.asdata(wr_address_i_int_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_0),
	.prn(vcc));
defparam \wraddress_b_bus[0] .is_wysiwyg = "true";
defparam \wraddress_b_bus[0] .power_up = "low";

dffeas \wraddress_b_bus[9] (
	.clk(clk),
	.d(ram_in_reg_1_1),
	.asdata(wr_address_i_int_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_9),
	.prn(vcc));
defparam \wraddress_b_bus[9] .is_wysiwyg = "true";
defparam \wraddress_b_bus[9] .power_up = "low";

dffeas \wraddress_b_bus[10] (
	.clk(clk),
	.d(ram_block6a0),
	.asdata(wr_address_i_int_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_10),
	.prn(vcc));
defparam \wraddress_b_bus[10] .is_wysiwyg = "true";
defparam \wraddress_b_bus[10] .power_up = "low";

dffeas \wraddress_b_bus[11] (
	.clk(clk),
	.d(ram_block6a1),
	.asdata(wr_address_i_int_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_11),
	.prn(vcc));
defparam \wraddress_b_bus[11] .is_wysiwyg = "true";
defparam \wraddress_b_bus[11] .power_up = "low";

dffeas \rdaddress_b_bus[0] (
	.clk(clk),
	.d(ram_in_reg_0_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_0),
	.prn(vcc));
defparam \rdaddress_b_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[0] .power_up = "low";

dffeas \rdaddress_b_bus[9] (
	.clk(clk),
	.d(ram_in_reg_1_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_9),
	.prn(vcc));
defparam \rdaddress_b_bus[9] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[9] .power_up = "low";

dffeas \rdaddress_b_bus[10] (
	.clk(clk),
	.d(ram_in_reg_2_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_10),
	.prn(vcc));
defparam \rdaddress_b_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[10] .power_up = "low";

dffeas \rdaddress_b_bus[11] (
	.clk(clk),
	.d(ram_in_reg_3_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_11),
	.prn(vcc));
defparam \rdaddress_b_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[11] .power_up = "low";

dffeas \a_ram_data_in_bus[46] (
	.clk(clk),
	.d(data_in_r_6),
	.asdata(ram_in_reg_6_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_46),
	.prn(vcc));
defparam \a_ram_data_in_bus[46] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[46] .power_up = "low";

dffeas \wraddress_a_bus[0] (
	.clk(clk),
	.d(wr_address_i_int_0),
	.asdata(ram_in_reg_0_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_0),
	.prn(vcc));
defparam \wraddress_a_bus[0] .is_wysiwyg = "true";
defparam \wraddress_a_bus[0] .power_up = "low";

dffeas \wraddress_a_bus[9] (
	.clk(clk),
	.d(wr_address_i_int_1),
	.asdata(ram_in_reg_1_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_9),
	.prn(vcc));
defparam \wraddress_a_bus[9] .is_wysiwyg = "true";
defparam \wraddress_a_bus[9] .power_up = "low";

dffeas \wraddress_a_bus[10] (
	.clk(clk),
	.d(wr_address_i_int_2),
	.asdata(ram_block6a0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_10),
	.prn(vcc));
defparam \wraddress_a_bus[10] .is_wysiwyg = "true";
defparam \wraddress_a_bus[10] .power_up = "low";

dffeas \wraddress_a_bus[11] (
	.clk(clk),
	.d(wr_address_i_int_3),
	.asdata(ram_block6a1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_11),
	.prn(vcc));
defparam \wraddress_a_bus[11] .is_wysiwyg = "true";
defparam \wraddress_a_bus[11] .power_up = "low";

dffeas \rdaddress_a_bus[0] (
	.clk(clk),
	.d(ram_in_reg_0_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_0),
	.prn(vcc));
defparam \rdaddress_a_bus[0] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[0] .power_up = "low";

dffeas \rdaddress_a_bus[9] (
	.clk(clk),
	.d(ram_in_reg_1_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_9),
	.prn(vcc));
defparam \rdaddress_a_bus[9] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[9] .power_up = "low";

dffeas \rdaddress_a_bus[10] (
	.clk(clk),
	.d(ram_in_reg_2_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_10),
	.prn(vcc));
defparam \rdaddress_a_bus[10] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[10] .power_up = "low";

dffeas \rdaddress_a_bus[11] (
	.clk(clk),
	.d(ram_in_reg_3_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_11),
	.prn(vcc));
defparam \rdaddress_a_bus[11] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[11] .power_up = "low";

dffeas \b_ram_data_in_bus[30] (
	.clk(clk),
	.d(ram_in_reg_6_2),
	.asdata(data_in_r_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_30),
	.prn(vcc));
defparam \b_ram_data_in_bus[30] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[30] .power_up = "low";

dffeas \wraddress_b_bus[12] (
	.clk(clk),
	.d(ram_in_reg_0_0),
	.asdata(wr_address_i_int_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_12),
	.prn(vcc));
defparam \wraddress_b_bus[12] .is_wysiwyg = "true";
defparam \wraddress_b_bus[12] .power_up = "low";

dffeas \wraddress_b_bus[5] (
	.clk(clk),
	.d(ram_in_reg_1_2),
	.asdata(wr_address_i_int_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_5),
	.prn(vcc));
defparam \wraddress_b_bus[5] .is_wysiwyg = "true";
defparam \wraddress_b_bus[5] .power_up = "low";

dffeas \rdaddress_b_bus[12] (
	.clk(clk),
	.d(ram_in_reg_0_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_12),
	.prn(vcc));
defparam \rdaddress_b_bus[12] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[12] .power_up = "low";

dffeas \rdaddress_b_bus[5] (
	.clk(clk),
	.d(ram_in_reg_1_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_5),
	.prn(vcc));
defparam \rdaddress_b_bus[5] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[5] .power_up = "low";

dffeas \a_ram_data_in_bus[30] (
	.clk(clk),
	.d(data_in_r_6),
	.asdata(ram_in_reg_6_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_30),
	.prn(vcc));
defparam \a_ram_data_in_bus[30] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[30] .power_up = "low";

dffeas \wraddress_a_bus[12] (
	.clk(clk),
	.d(wr_address_i_int_0),
	.asdata(ram_in_reg_0_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_12),
	.prn(vcc));
defparam \wraddress_a_bus[12] .is_wysiwyg = "true";
defparam \wraddress_a_bus[12] .power_up = "low";

dffeas \wraddress_a_bus[5] (
	.clk(clk),
	.d(wr_address_i_int_1),
	.asdata(ram_in_reg_1_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_5),
	.prn(vcc));
defparam \wraddress_a_bus[5] .is_wysiwyg = "true";
defparam \wraddress_a_bus[5] .power_up = "low";

dffeas \rdaddress_a_bus[12] (
	.clk(clk),
	.d(ram_in_reg_0_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_12),
	.prn(vcc));
defparam \rdaddress_a_bus[12] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[12] .power_up = "low";

dffeas \rdaddress_a_bus[5] (
	.clk(clk),
	.d(ram_in_reg_1_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_5),
	.prn(vcc));
defparam \rdaddress_a_bus[5] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[5] .power_up = "low";

dffeas \b_ram_data_in_bus[14] (
	.clk(clk),
	.d(ram_in_reg_6_3),
	.asdata(data_in_r_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_14),
	.prn(vcc));
defparam \b_ram_data_in_bus[14] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[14] .power_up = "low";

dffeas \wraddress_b_bus[1] (
	.clk(clk),
	.d(ram_in_reg_1_3),
	.asdata(wr_address_i_int_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_1),
	.prn(vcc));
defparam \wraddress_b_bus[1] .is_wysiwyg = "true";
defparam \wraddress_b_bus[1] .power_up = "low";

dffeas \rdaddress_b_bus[1] (
	.clk(clk),
	.d(ram_in_reg_1_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_1),
	.prn(vcc));
defparam \rdaddress_b_bus[1] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[1] .power_up = "low";

dffeas \a_ram_data_in_bus[14] (
	.clk(clk),
	.d(data_in_r_6),
	.asdata(ram_in_reg_6_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_14),
	.prn(vcc));
defparam \a_ram_data_in_bus[14] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[14] .power_up = "low";

dffeas \wraddress_a_bus[1] (
	.clk(clk),
	.d(wr_address_i_int_1),
	.asdata(ram_in_reg_1_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_1),
	.prn(vcc));
defparam \wraddress_a_bus[1] .is_wysiwyg = "true";
defparam \wraddress_a_bus[1] .power_up = "low";

dffeas \rdaddress_a_bus[1] (
	.clk(clk),
	.d(ram_in_reg_1_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_1),
	.prn(vcc));
defparam \rdaddress_a_bus[1] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[1] .power_up = "low";

dffeas \b_ram_data_in_bus[62] (
	.clk(clk),
	.d(ram_in_reg_6_0),
	.asdata(data_in_r_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_62),
	.prn(vcc));
defparam \b_ram_data_in_bus[62] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[62] .power_up = "low";

dffeas \wraddress_b_bus[13] (
	.clk(clk),
	.d(ram_in_reg_1_0),
	.asdata(wr_address_i_int_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_b_bus_13),
	.prn(vcc));
defparam \wraddress_b_bus[13] .is_wysiwyg = "true";
defparam \wraddress_b_bus[13] .power_up = "low";

dffeas \rdaddress_b_bus[13] (
	.clk(clk),
	.d(ram_in_reg_1_02),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_b_bus_13),
	.prn(vcc));
defparam \rdaddress_b_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_b_bus[13] .power_up = "low";

dffeas \a_ram_data_in_bus[62] (
	.clk(clk),
	.d(data_in_r_6),
	.asdata(ram_in_reg_6_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_62),
	.prn(vcc));
defparam \a_ram_data_in_bus[62] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[62] .power_up = "low";

dffeas \wraddress_a_bus[13] (
	.clk(clk),
	.d(wr_address_i_int_1),
	.asdata(ram_in_reg_1_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(wraddress_a_bus_13),
	.prn(vcc));
defparam \wraddress_a_bus[13] .is_wysiwyg = "true";
defparam \wraddress_a_bus[13] .power_up = "low";

dffeas \rdaddress_a_bus[13] (
	.clk(clk),
	.d(ram_in_reg_1_02),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(sel_anb_addr),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rdaddress_a_bus_13),
	.prn(vcc));
defparam \rdaddress_a_bus[13] .is_wysiwyg = "true";
defparam \rdaddress_a_bus[13] .power_up = "low";

dffeas \b_ram_data_in_bus[45] (
	.clk(clk),
	.d(ram_in_reg_5_1),
	.asdata(data_in_r_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_45),
	.prn(vcc));
defparam \b_ram_data_in_bus[45] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[45] .power_up = "low";

dffeas \a_ram_data_in_bus[45] (
	.clk(clk),
	.d(data_in_r_5),
	.asdata(ram_in_reg_5_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_45),
	.prn(vcc));
defparam \a_ram_data_in_bus[45] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[45] .power_up = "low";

dffeas \b_ram_data_in_bus[29] (
	.clk(clk),
	.d(ram_in_reg_5_2),
	.asdata(data_in_r_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_29),
	.prn(vcc));
defparam \b_ram_data_in_bus[29] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[29] .power_up = "low";

dffeas \a_ram_data_in_bus[29] (
	.clk(clk),
	.d(data_in_r_5),
	.asdata(ram_in_reg_5_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_29),
	.prn(vcc));
defparam \a_ram_data_in_bus[29] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[29] .power_up = "low";

dffeas \b_ram_data_in_bus[13] (
	.clk(clk),
	.d(ram_in_reg_5_3),
	.asdata(data_in_r_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_13),
	.prn(vcc));
defparam \b_ram_data_in_bus[13] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[13] .power_up = "low";

dffeas \a_ram_data_in_bus[13] (
	.clk(clk),
	.d(data_in_r_5),
	.asdata(ram_in_reg_5_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_13),
	.prn(vcc));
defparam \a_ram_data_in_bus[13] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[13] .power_up = "low";

dffeas \b_ram_data_in_bus[61] (
	.clk(clk),
	.d(ram_in_reg_5_0),
	.asdata(data_in_r_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_61),
	.prn(vcc));
defparam \b_ram_data_in_bus[61] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[61] .power_up = "low";

dffeas \a_ram_data_in_bus[61] (
	.clk(clk),
	.d(data_in_r_5),
	.asdata(ram_in_reg_5_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_61),
	.prn(vcc));
defparam \a_ram_data_in_bus[61] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[61] .power_up = "low";

dffeas \b_ram_data_in_bus[42] (
	.clk(clk),
	.d(ram_in_reg_2_1),
	.asdata(data_in_r_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_42),
	.prn(vcc));
defparam \b_ram_data_in_bus[42] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[42] .power_up = "low";

dffeas \a_ram_data_in_bus[42] (
	.clk(clk),
	.d(data_in_r_2),
	.asdata(ram_in_reg_2_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_42),
	.prn(vcc));
defparam \a_ram_data_in_bus[42] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[42] .power_up = "low";

dffeas \b_ram_data_in_bus[26] (
	.clk(clk),
	.d(ram_in_reg_2_2),
	.asdata(data_in_r_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_26),
	.prn(vcc));
defparam \b_ram_data_in_bus[26] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[26] .power_up = "low";

dffeas \a_ram_data_in_bus[26] (
	.clk(clk),
	.d(data_in_r_2),
	.asdata(ram_in_reg_2_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_26),
	.prn(vcc));
defparam \a_ram_data_in_bus[26] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[26] .power_up = "low";

dffeas \b_ram_data_in_bus[10] (
	.clk(clk),
	.d(ram_in_reg_2_3),
	.asdata(data_in_r_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_10),
	.prn(vcc));
defparam \b_ram_data_in_bus[10] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[10] .power_up = "low";

dffeas \a_ram_data_in_bus[10] (
	.clk(clk),
	.d(data_in_r_2),
	.asdata(ram_in_reg_2_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_10),
	.prn(vcc));
defparam \a_ram_data_in_bus[10] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[10] .power_up = "low";

dffeas \b_ram_data_in_bus[58] (
	.clk(clk),
	.d(ram_in_reg_2_0),
	.asdata(data_in_r_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_58),
	.prn(vcc));
defparam \b_ram_data_in_bus[58] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[58] .power_up = "low";

dffeas \a_ram_data_in_bus[58] (
	.clk(clk),
	.d(data_in_r_2),
	.asdata(ram_in_reg_2_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_58),
	.prn(vcc));
defparam \a_ram_data_in_bus[58] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[58] .power_up = "low";

dffeas \b_ram_data_in_bus[43] (
	.clk(clk),
	.d(ram_in_reg_3_1),
	.asdata(data_in_r_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_43),
	.prn(vcc));
defparam \b_ram_data_in_bus[43] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[43] .power_up = "low";

dffeas \a_ram_data_in_bus[43] (
	.clk(clk),
	.d(data_in_r_3),
	.asdata(ram_in_reg_3_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_43),
	.prn(vcc));
defparam \a_ram_data_in_bus[43] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[43] .power_up = "low";

dffeas \b_ram_data_in_bus[27] (
	.clk(clk),
	.d(ram_in_reg_3_2),
	.asdata(data_in_r_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_27),
	.prn(vcc));
defparam \b_ram_data_in_bus[27] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[27] .power_up = "low";

dffeas \a_ram_data_in_bus[27] (
	.clk(clk),
	.d(data_in_r_3),
	.asdata(ram_in_reg_3_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_27),
	.prn(vcc));
defparam \a_ram_data_in_bus[27] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[27] .power_up = "low";

dffeas \b_ram_data_in_bus[11] (
	.clk(clk),
	.d(ram_in_reg_3_3),
	.asdata(data_in_r_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_11),
	.prn(vcc));
defparam \b_ram_data_in_bus[11] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[11] .power_up = "low";

dffeas \a_ram_data_in_bus[11] (
	.clk(clk),
	.d(data_in_r_3),
	.asdata(ram_in_reg_3_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_11),
	.prn(vcc));
defparam \a_ram_data_in_bus[11] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[11] .power_up = "low";

dffeas \b_ram_data_in_bus[59] (
	.clk(clk),
	.d(ram_in_reg_3_0),
	.asdata(data_in_r_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_59),
	.prn(vcc));
defparam \b_ram_data_in_bus[59] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[59] .power_up = "low";

dffeas \a_ram_data_in_bus[59] (
	.clk(clk),
	.d(data_in_r_3),
	.asdata(ram_in_reg_3_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_59),
	.prn(vcc));
defparam \a_ram_data_in_bus[59] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[59] .power_up = "low";

dffeas \b_ram_data_in_bus[44] (
	.clk(clk),
	.d(ram_in_reg_4_1),
	.asdata(data_in_r_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_44),
	.prn(vcc));
defparam \b_ram_data_in_bus[44] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[44] .power_up = "low";

dffeas \a_ram_data_in_bus[44] (
	.clk(clk),
	.d(data_in_r_4),
	.asdata(ram_in_reg_4_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_44),
	.prn(vcc));
defparam \a_ram_data_in_bus[44] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[44] .power_up = "low";

dffeas \b_ram_data_in_bus[28] (
	.clk(clk),
	.d(ram_in_reg_4_2),
	.asdata(data_in_r_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_28),
	.prn(vcc));
defparam \b_ram_data_in_bus[28] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[28] .power_up = "low";

dffeas \a_ram_data_in_bus[28] (
	.clk(clk),
	.d(data_in_r_4),
	.asdata(ram_in_reg_4_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_28),
	.prn(vcc));
defparam \a_ram_data_in_bus[28] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[28] .power_up = "low";

dffeas \b_ram_data_in_bus[12] (
	.clk(clk),
	.d(ram_in_reg_4_3),
	.asdata(data_in_r_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_12),
	.prn(vcc));
defparam \b_ram_data_in_bus[12] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[12] .power_up = "low";

dffeas \a_ram_data_in_bus[12] (
	.clk(clk),
	.d(data_in_r_4),
	.asdata(ram_in_reg_4_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_12),
	.prn(vcc));
defparam \a_ram_data_in_bus[12] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[12] .power_up = "low";

dffeas \b_ram_data_in_bus[60] (
	.clk(clk),
	.d(ram_in_reg_4_0),
	.asdata(data_in_r_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_60),
	.prn(vcc));
defparam \b_ram_data_in_bus[60] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[60] .power_up = "low";

dffeas \a_ram_data_in_bus[60] (
	.clk(clk),
	.d(data_in_r_4),
	.asdata(ram_in_reg_4_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_60),
	.prn(vcc));
defparam \a_ram_data_in_bus[60] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[60] .power_up = "low";

dffeas \b_ram_data_in_bus[47] (
	.clk(clk),
	.d(ram_in_reg_7_1),
	.asdata(data_in_r_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_47),
	.prn(vcc));
defparam \b_ram_data_in_bus[47] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[47] .power_up = "low";

dffeas \a_ram_data_in_bus[47] (
	.clk(clk),
	.d(data_in_r_7),
	.asdata(ram_in_reg_7_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_47),
	.prn(vcc));
defparam \a_ram_data_in_bus[47] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[47] .power_up = "low";

dffeas \b_ram_data_in_bus[31] (
	.clk(clk),
	.d(ram_in_reg_7_2),
	.asdata(data_in_r_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_31),
	.prn(vcc));
defparam \b_ram_data_in_bus[31] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[31] .power_up = "low";

dffeas \a_ram_data_in_bus[31] (
	.clk(clk),
	.d(data_in_r_7),
	.asdata(ram_in_reg_7_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_31),
	.prn(vcc));
defparam \a_ram_data_in_bus[31] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[31] .power_up = "low";

dffeas \b_ram_data_in_bus[15] (
	.clk(clk),
	.d(ram_in_reg_7_3),
	.asdata(data_in_r_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_15),
	.prn(vcc));
defparam \b_ram_data_in_bus[15] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[15] .power_up = "low";

dffeas \a_ram_data_in_bus[15] (
	.clk(clk),
	.d(data_in_r_7),
	.asdata(ram_in_reg_7_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_15),
	.prn(vcc));
defparam \a_ram_data_in_bus[15] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[15] .power_up = "low";

dffeas \b_ram_data_in_bus[63] (
	.clk(clk),
	.d(ram_in_reg_7_0),
	.asdata(data_in_r_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_63),
	.prn(vcc));
defparam \b_ram_data_in_bus[63] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[63] .power_up = "low";

dffeas \a_ram_data_in_bus[63] (
	.clk(clk),
	.d(data_in_r_7),
	.asdata(ram_in_reg_7_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_63),
	.prn(vcc));
defparam \a_ram_data_in_bus[63] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[63] .power_up = "low";

dffeas \b_ram_data_in_bus[39] (
	.clk(clk),
	.d(ram_in_reg_7_5),
	.asdata(data_in_i_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_39),
	.prn(vcc));
defparam \b_ram_data_in_bus[39] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[39] .power_up = "low";

dffeas \a_ram_data_in_bus[39] (
	.clk(clk),
	.d(data_in_i_7),
	.asdata(ram_in_reg_7_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_39),
	.prn(vcc));
defparam \a_ram_data_in_bus[39] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[39] .power_up = "low";

dffeas \b_ram_data_in_bus[23] (
	.clk(clk),
	.d(ram_in_reg_7_6),
	.asdata(data_in_i_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_23),
	.prn(vcc));
defparam \b_ram_data_in_bus[23] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[23] .power_up = "low";

dffeas \a_ram_data_in_bus[23] (
	.clk(clk),
	.d(data_in_i_7),
	.asdata(ram_in_reg_7_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_23),
	.prn(vcc));
defparam \a_ram_data_in_bus[23] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[23] .power_up = "low";

dffeas \b_ram_data_in_bus[7] (
	.clk(clk),
	.d(ram_in_reg_7_7),
	.asdata(data_in_i_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_7),
	.prn(vcc));
defparam \b_ram_data_in_bus[7] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[7] .power_up = "low";

dffeas \a_ram_data_in_bus[7] (
	.clk(clk),
	.d(data_in_i_7),
	.asdata(ram_in_reg_7_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_7),
	.prn(vcc));
defparam \a_ram_data_in_bus[7] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[7] .power_up = "low";

dffeas \b_ram_data_in_bus[55] (
	.clk(clk),
	.d(ram_in_reg_7_4),
	.asdata(data_in_i_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_55),
	.prn(vcc));
defparam \b_ram_data_in_bus[55] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[55] .power_up = "low";

dffeas \a_ram_data_in_bus[55] (
	.clk(clk),
	.d(data_in_i_7),
	.asdata(ram_in_reg_7_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_55),
	.prn(vcc));
defparam \a_ram_data_in_bus[55] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[55] .power_up = "low";

dffeas \b_ram_data_in_bus[38] (
	.clk(clk),
	.d(ram_in_reg_6_5),
	.asdata(data_in_i_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_38),
	.prn(vcc));
defparam \b_ram_data_in_bus[38] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[38] .power_up = "low";

dffeas \a_ram_data_in_bus[38] (
	.clk(clk),
	.d(data_in_i_6),
	.asdata(ram_in_reg_6_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_38),
	.prn(vcc));
defparam \a_ram_data_in_bus[38] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[38] .power_up = "low";

dffeas \b_ram_data_in_bus[22] (
	.clk(clk),
	.d(ram_in_reg_6_6),
	.asdata(data_in_i_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_22),
	.prn(vcc));
defparam \b_ram_data_in_bus[22] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[22] .power_up = "low";

dffeas \a_ram_data_in_bus[22] (
	.clk(clk),
	.d(data_in_i_6),
	.asdata(ram_in_reg_6_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_22),
	.prn(vcc));
defparam \a_ram_data_in_bus[22] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[22] .power_up = "low";

dffeas \b_ram_data_in_bus[6] (
	.clk(clk),
	.d(ram_in_reg_6_7),
	.asdata(data_in_i_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_6),
	.prn(vcc));
defparam \b_ram_data_in_bus[6] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[6] .power_up = "low";

dffeas \a_ram_data_in_bus[6] (
	.clk(clk),
	.d(data_in_i_6),
	.asdata(ram_in_reg_6_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_6),
	.prn(vcc));
defparam \a_ram_data_in_bus[6] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[6] .power_up = "low";

dffeas \b_ram_data_in_bus[54] (
	.clk(clk),
	.d(ram_in_reg_6_4),
	.asdata(data_in_i_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_54),
	.prn(vcc));
defparam \b_ram_data_in_bus[54] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[54] .power_up = "low";

dffeas \a_ram_data_in_bus[54] (
	.clk(clk),
	.d(data_in_i_6),
	.asdata(ram_in_reg_6_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_54),
	.prn(vcc));
defparam \a_ram_data_in_bus[54] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[54] .power_up = "low";

dffeas \b_ram_data_in_bus[35] (
	.clk(clk),
	.d(ram_in_reg_3_5),
	.asdata(data_in_i_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_35),
	.prn(vcc));
defparam \b_ram_data_in_bus[35] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[35] .power_up = "low";

dffeas \a_ram_data_in_bus[35] (
	.clk(clk),
	.d(data_in_i_3),
	.asdata(ram_in_reg_3_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_35),
	.prn(vcc));
defparam \a_ram_data_in_bus[35] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[35] .power_up = "low";

dffeas \b_ram_data_in_bus[19] (
	.clk(clk),
	.d(ram_in_reg_3_6),
	.asdata(data_in_i_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_19),
	.prn(vcc));
defparam \b_ram_data_in_bus[19] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[19] .power_up = "low";

dffeas \a_ram_data_in_bus[19] (
	.clk(clk),
	.d(data_in_i_3),
	.asdata(ram_in_reg_3_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_19),
	.prn(vcc));
defparam \a_ram_data_in_bus[19] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[19] .power_up = "low";

dffeas \b_ram_data_in_bus[3] (
	.clk(clk),
	.d(ram_in_reg_3_7),
	.asdata(data_in_i_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_3),
	.prn(vcc));
defparam \b_ram_data_in_bus[3] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[3] .power_up = "low";

dffeas \a_ram_data_in_bus[3] (
	.clk(clk),
	.d(data_in_i_3),
	.asdata(ram_in_reg_3_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_3),
	.prn(vcc));
defparam \a_ram_data_in_bus[3] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[3] .power_up = "low";

dffeas \b_ram_data_in_bus[51] (
	.clk(clk),
	.d(ram_in_reg_3_4),
	.asdata(data_in_i_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_51),
	.prn(vcc));
defparam \b_ram_data_in_bus[51] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[51] .power_up = "low";

dffeas \a_ram_data_in_bus[51] (
	.clk(clk),
	.d(data_in_i_3),
	.asdata(ram_in_reg_3_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_51),
	.prn(vcc));
defparam \a_ram_data_in_bus[51] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[51] .power_up = "low";

dffeas \b_ram_data_in_bus[36] (
	.clk(clk),
	.d(ram_in_reg_4_5),
	.asdata(data_in_i_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_36),
	.prn(vcc));
defparam \b_ram_data_in_bus[36] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[36] .power_up = "low";

dffeas \a_ram_data_in_bus[36] (
	.clk(clk),
	.d(data_in_i_4),
	.asdata(ram_in_reg_4_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_36),
	.prn(vcc));
defparam \a_ram_data_in_bus[36] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[36] .power_up = "low";

dffeas \b_ram_data_in_bus[20] (
	.clk(clk),
	.d(ram_in_reg_4_6),
	.asdata(data_in_i_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_20),
	.prn(vcc));
defparam \b_ram_data_in_bus[20] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[20] .power_up = "low";

dffeas \a_ram_data_in_bus[20] (
	.clk(clk),
	.d(data_in_i_4),
	.asdata(ram_in_reg_4_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_20),
	.prn(vcc));
defparam \a_ram_data_in_bus[20] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[20] .power_up = "low";

dffeas \b_ram_data_in_bus[4] (
	.clk(clk),
	.d(ram_in_reg_4_7),
	.asdata(data_in_i_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_4),
	.prn(vcc));
defparam \b_ram_data_in_bus[4] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[4] .power_up = "low";

dffeas \a_ram_data_in_bus[4] (
	.clk(clk),
	.d(data_in_i_4),
	.asdata(ram_in_reg_4_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_4),
	.prn(vcc));
defparam \a_ram_data_in_bus[4] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[4] .power_up = "low";

dffeas \b_ram_data_in_bus[52] (
	.clk(clk),
	.d(ram_in_reg_4_4),
	.asdata(data_in_i_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_52),
	.prn(vcc));
defparam \b_ram_data_in_bus[52] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[52] .power_up = "low";

dffeas \a_ram_data_in_bus[52] (
	.clk(clk),
	.d(data_in_i_4),
	.asdata(ram_in_reg_4_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_52),
	.prn(vcc));
defparam \a_ram_data_in_bus[52] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[52] .power_up = "low";

dffeas \b_ram_data_in_bus[37] (
	.clk(clk),
	.d(ram_in_reg_5_5),
	.asdata(data_in_i_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_37),
	.prn(vcc));
defparam \b_ram_data_in_bus[37] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[37] .power_up = "low";

dffeas \a_ram_data_in_bus[37] (
	.clk(clk),
	.d(data_in_i_5),
	.asdata(ram_in_reg_5_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_37),
	.prn(vcc));
defparam \a_ram_data_in_bus[37] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[37] .power_up = "low";

dffeas \b_ram_data_in_bus[21] (
	.clk(clk),
	.d(ram_in_reg_5_6),
	.asdata(data_in_i_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_21),
	.prn(vcc));
defparam \b_ram_data_in_bus[21] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[21] .power_up = "low";

dffeas \a_ram_data_in_bus[21] (
	.clk(clk),
	.d(data_in_i_5),
	.asdata(ram_in_reg_5_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_21),
	.prn(vcc));
defparam \a_ram_data_in_bus[21] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[21] .power_up = "low";

dffeas \b_ram_data_in_bus[5] (
	.clk(clk),
	.d(ram_in_reg_5_7),
	.asdata(data_in_i_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_5),
	.prn(vcc));
defparam \b_ram_data_in_bus[5] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[5] .power_up = "low";

dffeas \a_ram_data_in_bus[5] (
	.clk(clk),
	.d(data_in_i_5),
	.asdata(ram_in_reg_5_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_5),
	.prn(vcc));
defparam \a_ram_data_in_bus[5] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[5] .power_up = "low";

dffeas \b_ram_data_in_bus[53] (
	.clk(clk),
	.d(ram_in_reg_5_4),
	.asdata(data_in_i_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_53),
	.prn(vcc));
defparam \b_ram_data_in_bus[53] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[53] .power_up = "low";

dffeas \a_ram_data_in_bus[53] (
	.clk(clk),
	.d(data_in_i_5),
	.asdata(ram_in_reg_5_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_53),
	.prn(vcc));
defparam \a_ram_data_in_bus[53] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[53] .power_up = "low";

dffeas \b_ram_data_in_bus[34] (
	.clk(clk),
	.d(ram_in_reg_2_5),
	.asdata(data_in_i_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_34),
	.prn(vcc));
defparam \b_ram_data_in_bus[34] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[34] .power_up = "low";

dffeas \a_ram_data_in_bus[34] (
	.clk(clk),
	.d(data_in_i_2),
	.asdata(ram_in_reg_2_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_34),
	.prn(vcc));
defparam \a_ram_data_in_bus[34] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[34] .power_up = "low";

dffeas \b_ram_data_in_bus[18] (
	.clk(clk),
	.d(ram_in_reg_2_6),
	.asdata(data_in_i_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_18),
	.prn(vcc));
defparam \b_ram_data_in_bus[18] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[18] .power_up = "low";

dffeas \a_ram_data_in_bus[18] (
	.clk(clk),
	.d(data_in_i_2),
	.asdata(ram_in_reg_2_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_18),
	.prn(vcc));
defparam \a_ram_data_in_bus[18] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[18] .power_up = "low";

dffeas \b_ram_data_in_bus[2] (
	.clk(clk),
	.d(ram_in_reg_2_7),
	.asdata(data_in_i_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_2),
	.prn(vcc));
defparam \b_ram_data_in_bus[2] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[2] .power_up = "low";

dffeas \a_ram_data_in_bus[2] (
	.clk(clk),
	.d(data_in_i_2),
	.asdata(ram_in_reg_2_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_2),
	.prn(vcc));
defparam \a_ram_data_in_bus[2] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[2] .power_up = "low";

dffeas \b_ram_data_in_bus[50] (
	.clk(clk),
	.d(ram_in_reg_2_4),
	.asdata(data_in_i_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_50),
	.prn(vcc));
defparam \b_ram_data_in_bus[50] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[50] .power_up = "low";

dffeas \a_ram_data_in_bus[50] (
	.clk(clk),
	.d(data_in_i_2),
	.asdata(ram_in_reg_2_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_50),
	.prn(vcc));
defparam \a_ram_data_in_bus[50] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[50] .power_up = "low";

dffeas \b_ram_data_in_bus[24] (
	.clk(clk),
	.d(ram_in_reg_0_2),
	.asdata(data_in_r_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_24),
	.prn(vcc));
defparam \b_ram_data_in_bus[24] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[24] .power_up = "low";

dffeas \a_ram_data_in_bus[24] (
	.clk(clk),
	.d(data_in_r_0),
	.asdata(ram_in_reg_0_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_24),
	.prn(vcc));
defparam \a_ram_data_in_bus[24] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[24] .power_up = "low";

dffeas \b_ram_data_in_bus[8] (
	.clk(clk),
	.d(ram_in_reg_0_3),
	.asdata(data_in_r_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_8),
	.prn(vcc));
defparam \b_ram_data_in_bus[8] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[8] .power_up = "low";

dffeas \a_ram_data_in_bus[8] (
	.clk(clk),
	.d(data_in_r_0),
	.asdata(ram_in_reg_0_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_8),
	.prn(vcc));
defparam \a_ram_data_in_bus[8] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[8] .power_up = "low";

dffeas \b_ram_data_in_bus[56] (
	.clk(clk),
	.d(ram_in_reg_0_02),
	.asdata(data_in_r_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_56),
	.prn(vcc));
defparam \b_ram_data_in_bus[56] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[56] .power_up = "low";

dffeas \a_ram_data_in_bus[56] (
	.clk(clk),
	.d(data_in_r_0),
	.asdata(ram_in_reg_0_02),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_56),
	.prn(vcc));
defparam \a_ram_data_in_bus[56] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[56] .power_up = "low";

dffeas \b_ram_data_in_bus[40] (
	.clk(clk),
	.d(ram_in_reg_0_12),
	.asdata(data_in_r_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_40),
	.prn(vcc));
defparam \b_ram_data_in_bus[40] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[40] .power_up = "low";

dffeas \a_ram_data_in_bus[40] (
	.clk(clk),
	.d(data_in_r_0),
	.asdata(ram_in_reg_0_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_40),
	.prn(vcc));
defparam \a_ram_data_in_bus[40] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[40] .power_up = "low";

dffeas \b_ram_data_in_bus[25] (
	.clk(clk),
	.d(ram_in_reg_1_21),
	.asdata(data_in_r_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_25),
	.prn(vcc));
defparam \b_ram_data_in_bus[25] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[25] .power_up = "low";

dffeas \a_ram_data_in_bus[25] (
	.clk(clk),
	.d(data_in_r_1),
	.asdata(ram_in_reg_1_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_25),
	.prn(vcc));
defparam \a_ram_data_in_bus[25] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[25] .power_up = "low";

dffeas \b_ram_data_in_bus[9] (
	.clk(clk),
	.d(ram_in_reg_1_31),
	.asdata(data_in_r_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_9),
	.prn(vcc));
defparam \b_ram_data_in_bus[9] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[9] .power_up = "low";

dffeas \a_ram_data_in_bus[9] (
	.clk(clk),
	.d(data_in_r_1),
	.asdata(ram_in_reg_1_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_9),
	.prn(vcc));
defparam \a_ram_data_in_bus[9] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[9] .power_up = "low";

dffeas \b_ram_data_in_bus[57] (
	.clk(clk),
	.d(ram_in_reg_1_01),
	.asdata(data_in_r_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_57),
	.prn(vcc));
defparam \b_ram_data_in_bus[57] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[57] .power_up = "low";

dffeas \a_ram_data_in_bus[57] (
	.clk(clk),
	.d(data_in_r_1),
	.asdata(ram_in_reg_1_01),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_57),
	.prn(vcc));
defparam \a_ram_data_in_bus[57] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[57] .power_up = "low";

dffeas \b_ram_data_in_bus[41] (
	.clk(clk),
	.d(ram_in_reg_1_11),
	.asdata(data_in_r_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_41),
	.prn(vcc));
defparam \b_ram_data_in_bus[41] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[41] .power_up = "low";

dffeas \a_ram_data_in_bus[41] (
	.clk(clk),
	.d(data_in_r_1),
	.asdata(ram_in_reg_1_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_41),
	.prn(vcc));
defparam \a_ram_data_in_bus[41] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[41] .power_up = "low";

dffeas \b_ram_data_in_bus[0] (
	.clk(clk),
	.d(ram_in_reg_0_7),
	.asdata(data_in_i_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_0),
	.prn(vcc));
defparam \b_ram_data_in_bus[0] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[0] .power_up = "low";

dffeas \a_ram_data_in_bus[0] (
	.clk(clk),
	.d(data_in_i_0),
	.asdata(ram_in_reg_0_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_0),
	.prn(vcc));
defparam \a_ram_data_in_bus[0] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[0] .power_up = "low";

dffeas \b_ram_data_in_bus[48] (
	.clk(clk),
	.d(ram_in_reg_0_4),
	.asdata(data_in_i_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_48),
	.prn(vcc));
defparam \b_ram_data_in_bus[48] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[48] .power_up = "low";

dffeas \a_ram_data_in_bus[48] (
	.clk(clk),
	.d(data_in_i_0),
	.asdata(ram_in_reg_0_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_48),
	.prn(vcc));
defparam \a_ram_data_in_bus[48] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[48] .power_up = "low";

dffeas \b_ram_data_in_bus[32] (
	.clk(clk),
	.d(ram_in_reg_0_5),
	.asdata(data_in_i_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_32),
	.prn(vcc));
defparam \b_ram_data_in_bus[32] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[32] .power_up = "low";

dffeas \a_ram_data_in_bus[32] (
	.clk(clk),
	.d(data_in_i_0),
	.asdata(ram_in_reg_0_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_32),
	.prn(vcc));
defparam \a_ram_data_in_bus[32] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[32] .power_up = "low";

dffeas \b_ram_data_in_bus[16] (
	.clk(clk),
	.d(ram_in_reg_0_6),
	.asdata(data_in_i_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_16),
	.prn(vcc));
defparam \b_ram_data_in_bus[16] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[16] .power_up = "low";

dffeas \a_ram_data_in_bus[16] (
	.clk(clk),
	.d(data_in_i_0),
	.asdata(ram_in_reg_0_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_16),
	.prn(vcc));
defparam \a_ram_data_in_bus[16] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[16] .power_up = "low";

dffeas \b_ram_data_in_bus[1] (
	.clk(clk),
	.d(ram_in_reg_1_7),
	.asdata(data_in_i_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_1),
	.prn(vcc));
defparam \b_ram_data_in_bus[1] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[1] .power_up = "low";

dffeas \a_ram_data_in_bus[1] (
	.clk(clk),
	.d(data_in_i_1),
	.asdata(ram_in_reg_1_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_1),
	.prn(vcc));
defparam \a_ram_data_in_bus[1] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[1] .power_up = "low";

dffeas \b_ram_data_in_bus[49] (
	.clk(clk),
	.d(ram_in_reg_1_4),
	.asdata(data_in_i_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_49),
	.prn(vcc));
defparam \b_ram_data_in_bus[49] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[49] .power_up = "low";

dffeas \a_ram_data_in_bus[49] (
	.clk(clk),
	.d(data_in_i_1),
	.asdata(ram_in_reg_1_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_49),
	.prn(vcc));
defparam \a_ram_data_in_bus[49] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[49] .power_up = "low";

dffeas \b_ram_data_in_bus[33] (
	.clk(clk),
	.d(ram_in_reg_1_5),
	.asdata(data_in_i_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_33),
	.prn(vcc));
defparam \b_ram_data_in_bus[33] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[33] .power_up = "low";

dffeas \a_ram_data_in_bus[33] (
	.clk(clk),
	.d(data_in_i_1),
	.asdata(ram_in_reg_1_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_33),
	.prn(vcc));
defparam \a_ram_data_in_bus[33] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[33] .power_up = "low";

dffeas \b_ram_data_in_bus[17] (
	.clk(clk),
	.d(ram_in_reg_1_6),
	.asdata(data_in_i_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(b_ram_data_in_bus_17),
	.prn(vcc));
defparam \b_ram_data_in_bus[17] .is_wysiwyg = "true";
defparam \b_ram_data_in_bus[17] .power_up = "low";

dffeas \a_ram_data_in_bus[17] (
	.clk(clk),
	.d(data_in_i_1),
	.asdata(ram_in_reg_1_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!ram_a_not_b_vec_1),
	.ena(!global_clock_enable),
	.q(a_ram_data_in_bus_17),
	.prn(vcc));
defparam \a_ram_data_in_bus[17] .is_wysiwyg = "true";
defparam \a_ram_data_in_bus[17] .power_up = "low";

dffeas \ram_data_out1[14] (
	.clk(clk),
	.d(\ram_data_out1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_14),
	.prn(vcc));
defparam \ram_data_out1[14] .is_wysiwyg = "true";
defparam \ram_data_out1[14] .power_up = "low";

dffeas \ram_data_out2[14] (
	.clk(clk),
	.d(\ram_data_out2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_14),
	.prn(vcc));
defparam \ram_data_out2[14] .is_wysiwyg = "true";
defparam \ram_data_out2[14] .power_up = "low";

dffeas \ram_data_out3[14] (
	.clk(clk),
	.d(\ram_data_out3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_14),
	.prn(vcc));
defparam \ram_data_out3[14] .is_wysiwyg = "true";
defparam \ram_data_out3[14] .power_up = "low";

dffeas \ram_data_out0[14] (
	.clk(clk),
	.d(\ram_data_out0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_14),
	.prn(vcc));
defparam \ram_data_out0[14] .is_wysiwyg = "true";
defparam \ram_data_out0[14] .power_up = "low";

dffeas \ram_data_out1[13] (
	.clk(clk),
	.d(\ram_data_out1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_13),
	.prn(vcc));
defparam \ram_data_out1[13] .is_wysiwyg = "true";
defparam \ram_data_out1[13] .power_up = "low";

dffeas \ram_data_out2[13] (
	.clk(clk),
	.d(\ram_data_out2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_13),
	.prn(vcc));
defparam \ram_data_out2[13] .is_wysiwyg = "true";
defparam \ram_data_out2[13] .power_up = "low";

dffeas \ram_data_out3[13] (
	.clk(clk),
	.d(\ram_data_out3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_13),
	.prn(vcc));
defparam \ram_data_out3[13] .is_wysiwyg = "true";
defparam \ram_data_out3[13] .power_up = "low";

dffeas \ram_data_out0[13] (
	.clk(clk),
	.d(\ram_data_out0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_13),
	.prn(vcc));
defparam \ram_data_out0[13] .is_wysiwyg = "true";
defparam \ram_data_out0[13] .power_up = "low";

dffeas \ram_data_out1[10] (
	.clk(clk),
	.d(\ram_data_out1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_10),
	.prn(vcc));
defparam \ram_data_out1[10] .is_wysiwyg = "true";
defparam \ram_data_out1[10] .power_up = "low";

dffeas \ram_data_out2[10] (
	.clk(clk),
	.d(\ram_data_out2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_10),
	.prn(vcc));
defparam \ram_data_out2[10] .is_wysiwyg = "true";
defparam \ram_data_out2[10] .power_up = "low";

dffeas \ram_data_out3[10] (
	.clk(clk),
	.d(\ram_data_out3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_10),
	.prn(vcc));
defparam \ram_data_out3[10] .is_wysiwyg = "true";
defparam \ram_data_out3[10] .power_up = "low";

dffeas \ram_data_out0[10] (
	.clk(clk),
	.d(\ram_data_out0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_10),
	.prn(vcc));
defparam \ram_data_out0[10] .is_wysiwyg = "true";
defparam \ram_data_out0[10] .power_up = "low";

dffeas \ram_data_out1[11] (
	.clk(clk),
	.d(\ram_data_out1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_11),
	.prn(vcc));
defparam \ram_data_out1[11] .is_wysiwyg = "true";
defparam \ram_data_out1[11] .power_up = "low";

dffeas \ram_data_out2[11] (
	.clk(clk),
	.d(\ram_data_out2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_11),
	.prn(vcc));
defparam \ram_data_out2[11] .is_wysiwyg = "true";
defparam \ram_data_out2[11] .power_up = "low";

dffeas \ram_data_out3[11] (
	.clk(clk),
	.d(\ram_data_out3~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_11),
	.prn(vcc));
defparam \ram_data_out3[11] .is_wysiwyg = "true";
defparam \ram_data_out3[11] .power_up = "low";

dffeas \ram_data_out0[11] (
	.clk(clk),
	.d(\ram_data_out0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_11),
	.prn(vcc));
defparam \ram_data_out0[11] .is_wysiwyg = "true";
defparam \ram_data_out0[11] .power_up = "low";

dffeas \ram_data_out1[12] (
	.clk(clk),
	.d(\ram_data_out1~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_12),
	.prn(vcc));
defparam \ram_data_out1[12] .is_wysiwyg = "true";
defparam \ram_data_out1[12] .power_up = "low";

dffeas \ram_data_out2[12] (
	.clk(clk),
	.d(\ram_data_out2~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_12),
	.prn(vcc));
defparam \ram_data_out2[12] .is_wysiwyg = "true";
defparam \ram_data_out2[12] .power_up = "low";

dffeas \ram_data_out3[12] (
	.clk(clk),
	.d(\ram_data_out3~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_12),
	.prn(vcc));
defparam \ram_data_out3[12] .is_wysiwyg = "true";
defparam \ram_data_out3[12] .power_up = "low";

dffeas \ram_data_out0[12] (
	.clk(clk),
	.d(\ram_data_out0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_12),
	.prn(vcc));
defparam \ram_data_out0[12] .is_wysiwyg = "true";
defparam \ram_data_out0[12] .power_up = "low";

dffeas \ram_data_out1[15] (
	.clk(clk),
	.d(\ram_data_out1~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_15),
	.prn(vcc));
defparam \ram_data_out1[15] .is_wysiwyg = "true";
defparam \ram_data_out1[15] .power_up = "low";

dffeas \ram_data_out2[15] (
	.clk(clk),
	.d(\ram_data_out2~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_15),
	.prn(vcc));
defparam \ram_data_out2[15] .is_wysiwyg = "true";
defparam \ram_data_out2[15] .power_up = "low";

dffeas \ram_data_out3[15] (
	.clk(clk),
	.d(\ram_data_out3~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_15),
	.prn(vcc));
defparam \ram_data_out3[15] .is_wysiwyg = "true";
defparam \ram_data_out3[15] .power_up = "low";

dffeas \ram_data_out0[15] (
	.clk(clk),
	.d(\ram_data_out0~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_15),
	.prn(vcc));
defparam \ram_data_out0[15] .is_wysiwyg = "true";
defparam \ram_data_out0[15] .power_up = "low";

dffeas \ram_data_out1[7] (
	.clk(clk),
	.d(\ram_data_out1~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_7),
	.prn(vcc));
defparam \ram_data_out1[7] .is_wysiwyg = "true";
defparam \ram_data_out1[7] .power_up = "low";

dffeas \ram_data_out2[7] (
	.clk(clk),
	.d(\ram_data_out2~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_7),
	.prn(vcc));
defparam \ram_data_out2[7] .is_wysiwyg = "true";
defparam \ram_data_out2[7] .power_up = "low";

dffeas \ram_data_out3[7] (
	.clk(clk),
	.d(\ram_data_out3~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_7),
	.prn(vcc));
defparam \ram_data_out3[7] .is_wysiwyg = "true";
defparam \ram_data_out3[7] .power_up = "low";

dffeas \ram_data_out0[7] (
	.clk(clk),
	.d(\ram_data_out0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_7),
	.prn(vcc));
defparam \ram_data_out0[7] .is_wysiwyg = "true";
defparam \ram_data_out0[7] .power_up = "low";

dffeas \ram_data_out1[6] (
	.clk(clk),
	.d(\ram_data_out1~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_6),
	.prn(vcc));
defparam \ram_data_out1[6] .is_wysiwyg = "true";
defparam \ram_data_out1[6] .power_up = "low";

dffeas \ram_data_out2[6] (
	.clk(clk),
	.d(\ram_data_out2~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_6),
	.prn(vcc));
defparam \ram_data_out2[6] .is_wysiwyg = "true";
defparam \ram_data_out2[6] .power_up = "low";

dffeas \ram_data_out3[6] (
	.clk(clk),
	.d(\ram_data_out3~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_6),
	.prn(vcc));
defparam \ram_data_out3[6] .is_wysiwyg = "true";
defparam \ram_data_out3[6] .power_up = "low";

dffeas \ram_data_out0[6] (
	.clk(clk),
	.d(\ram_data_out0~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_6),
	.prn(vcc));
defparam \ram_data_out0[6] .is_wysiwyg = "true";
defparam \ram_data_out0[6] .power_up = "low";

dffeas \ram_data_out1[3] (
	.clk(clk),
	.d(\ram_data_out1~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_3),
	.prn(vcc));
defparam \ram_data_out1[3] .is_wysiwyg = "true";
defparam \ram_data_out1[3] .power_up = "low";

dffeas \ram_data_out2[3] (
	.clk(clk),
	.d(\ram_data_out2~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_3),
	.prn(vcc));
defparam \ram_data_out2[3] .is_wysiwyg = "true";
defparam \ram_data_out2[3] .power_up = "low";

dffeas \ram_data_out3[3] (
	.clk(clk),
	.d(\ram_data_out3~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_3),
	.prn(vcc));
defparam \ram_data_out3[3] .is_wysiwyg = "true";
defparam \ram_data_out3[3] .power_up = "low";

dffeas \ram_data_out0[3] (
	.clk(clk),
	.d(\ram_data_out0~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_3),
	.prn(vcc));
defparam \ram_data_out0[3] .is_wysiwyg = "true";
defparam \ram_data_out0[3] .power_up = "low";

dffeas \ram_data_out1[4] (
	.clk(clk),
	.d(\ram_data_out1~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_4),
	.prn(vcc));
defparam \ram_data_out1[4] .is_wysiwyg = "true";
defparam \ram_data_out1[4] .power_up = "low";

dffeas \ram_data_out2[4] (
	.clk(clk),
	.d(\ram_data_out2~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_4),
	.prn(vcc));
defparam \ram_data_out2[4] .is_wysiwyg = "true";
defparam \ram_data_out2[4] .power_up = "low";

dffeas \ram_data_out3[4] (
	.clk(clk),
	.d(\ram_data_out3~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_4),
	.prn(vcc));
defparam \ram_data_out3[4] .is_wysiwyg = "true";
defparam \ram_data_out3[4] .power_up = "low";

dffeas \ram_data_out0[4] (
	.clk(clk),
	.d(\ram_data_out0~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_4),
	.prn(vcc));
defparam \ram_data_out0[4] .is_wysiwyg = "true";
defparam \ram_data_out0[4] .power_up = "low";

dffeas \ram_data_out1[5] (
	.clk(clk),
	.d(\ram_data_out1~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_5),
	.prn(vcc));
defparam \ram_data_out1[5] .is_wysiwyg = "true";
defparam \ram_data_out1[5] .power_up = "low";

dffeas \ram_data_out2[5] (
	.clk(clk),
	.d(\ram_data_out2~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_5),
	.prn(vcc));
defparam \ram_data_out2[5] .is_wysiwyg = "true";
defparam \ram_data_out2[5] .power_up = "low";

dffeas \ram_data_out3[5] (
	.clk(clk),
	.d(\ram_data_out3~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_5),
	.prn(vcc));
defparam \ram_data_out3[5] .is_wysiwyg = "true";
defparam \ram_data_out3[5] .power_up = "low";

dffeas \ram_data_out0[5] (
	.clk(clk),
	.d(\ram_data_out0~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_5),
	.prn(vcc));
defparam \ram_data_out0[5] .is_wysiwyg = "true";
defparam \ram_data_out0[5] .power_up = "low";

dffeas \ram_data_out1[2] (
	.clk(clk),
	.d(\ram_data_out1~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_2),
	.prn(vcc));
defparam \ram_data_out1[2] .is_wysiwyg = "true";
defparam \ram_data_out1[2] .power_up = "low";

dffeas \ram_data_out2[2] (
	.clk(clk),
	.d(\ram_data_out2~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_2),
	.prn(vcc));
defparam \ram_data_out2[2] .is_wysiwyg = "true";
defparam \ram_data_out2[2] .power_up = "low";

dffeas \ram_data_out3[2] (
	.clk(clk),
	.d(\ram_data_out3~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_2),
	.prn(vcc));
defparam \ram_data_out3[2] .is_wysiwyg = "true";
defparam \ram_data_out3[2] .power_up = "low";

dffeas \ram_data_out0[2] (
	.clk(clk),
	.d(\ram_data_out0~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_2),
	.prn(vcc));
defparam \ram_data_out0[2] .is_wysiwyg = "true";
defparam \ram_data_out0[2] .power_up = "low";

dffeas \ram_data_out2[8] (
	.clk(clk),
	.d(\ram_data_out2~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_8),
	.prn(vcc));
defparam \ram_data_out2[8] .is_wysiwyg = "true";
defparam \ram_data_out2[8] .power_up = "low";

dffeas \ram_data_out3[8] (
	.clk(clk),
	.d(\ram_data_out3~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_8),
	.prn(vcc));
defparam \ram_data_out3[8] .is_wysiwyg = "true";
defparam \ram_data_out3[8] .power_up = "low";

dffeas \ram_data_out0[8] (
	.clk(clk),
	.d(\ram_data_out0~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_8),
	.prn(vcc));
defparam \ram_data_out0[8] .is_wysiwyg = "true";
defparam \ram_data_out0[8] .power_up = "low";

dffeas \ram_data_out1[8] (
	.clk(clk),
	.d(\ram_data_out1~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_8),
	.prn(vcc));
defparam \ram_data_out1[8] .is_wysiwyg = "true";
defparam \ram_data_out1[8] .power_up = "low";

dffeas \ram_data_out2[9] (
	.clk(clk),
	.d(\ram_data_out2~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_9),
	.prn(vcc));
defparam \ram_data_out2[9] .is_wysiwyg = "true";
defparam \ram_data_out2[9] .power_up = "low";

dffeas \ram_data_out3[9] (
	.clk(clk),
	.d(\ram_data_out3~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_9),
	.prn(vcc));
defparam \ram_data_out3[9] .is_wysiwyg = "true";
defparam \ram_data_out3[9] .power_up = "low";

dffeas \ram_data_out0[9] (
	.clk(clk),
	.d(\ram_data_out0~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_9),
	.prn(vcc));
defparam \ram_data_out0[9] .is_wysiwyg = "true";
defparam \ram_data_out0[9] .power_up = "low";

dffeas \ram_data_out1[9] (
	.clk(clk),
	.d(\ram_data_out1~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_9),
	.prn(vcc));
defparam \ram_data_out1[9] .is_wysiwyg = "true";
defparam \ram_data_out1[9] .power_up = "low";

dffeas \ram_data_out3[0] (
	.clk(clk),
	.d(\ram_data_out3~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_0),
	.prn(vcc));
defparam \ram_data_out3[0] .is_wysiwyg = "true";
defparam \ram_data_out3[0] .power_up = "low";

dffeas \ram_data_out0[0] (
	.clk(clk),
	.d(\ram_data_out0~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_0),
	.prn(vcc));
defparam \ram_data_out0[0] .is_wysiwyg = "true";
defparam \ram_data_out0[0] .power_up = "low";

dffeas \ram_data_out1[0] (
	.clk(clk),
	.d(\ram_data_out1~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_0),
	.prn(vcc));
defparam \ram_data_out1[0] .is_wysiwyg = "true";
defparam \ram_data_out1[0] .power_up = "low";

dffeas \ram_data_out2[0] (
	.clk(clk),
	.d(\ram_data_out2~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_0),
	.prn(vcc));
defparam \ram_data_out2[0] .is_wysiwyg = "true";
defparam \ram_data_out2[0] .power_up = "low";

dffeas \ram_data_out3[1] (
	.clk(clk),
	.d(\ram_data_out3~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out3_1),
	.prn(vcc));
defparam \ram_data_out3[1] .is_wysiwyg = "true";
defparam \ram_data_out3[1] .power_up = "low";

dffeas \ram_data_out0[1] (
	.clk(clk),
	.d(\ram_data_out0~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out0_1),
	.prn(vcc));
defparam \ram_data_out0[1] .is_wysiwyg = "true";
defparam \ram_data_out0[1] .power_up = "low";

dffeas \ram_data_out1[1] (
	.clk(clk),
	.d(\ram_data_out1~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out1_1),
	.prn(vcc));
defparam \ram_data_out1[1] .is_wysiwyg = "true";
defparam \ram_data_out1[1] .power_up = "low";

dffeas \ram_data_out2[1] (
	.clk(clk),
	.d(\ram_data_out2~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_data_out2_1),
	.prn(vcc));
defparam \ram_data_out2[1] .is_wysiwyg = "true";
defparam \ram_data_out2[1] .power_up = "low";

cyclonev_lcell_comb \ram_data_out1~0 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_14),
	.datad(!q_b_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~0 .extended_lut = "off";
defparam \ram_data_out1~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~0 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~0 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_142),
	.datad(!q_b_143),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~0 .extended_lut = "off";
defparam \ram_data_out2~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~0 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~0 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_144),
	.datad(!q_b_145),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~0 .extended_lut = "off";
defparam \ram_data_out3~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~0 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~0 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_146),
	.datad(!q_b_147),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~0 .extended_lut = "off";
defparam \ram_data_out0~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~0 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~1 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_13),
	.datad(!q_b_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~1 .extended_lut = "off";
defparam \ram_data_out1~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~1 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~1 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_132),
	.datad(!q_b_133),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~1 .extended_lut = "off";
defparam \ram_data_out2~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~1 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~1 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_134),
	.datad(!q_b_135),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~1 .extended_lut = "off";
defparam \ram_data_out3~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~1 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~1 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_136),
	.datad(!q_b_137),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~1 .extended_lut = "off";
defparam \ram_data_out0~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~1 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~2 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_10),
	.datad(!q_b_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~2 .extended_lut = "off";
defparam \ram_data_out1~2 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~2 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~2 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_102),
	.datad(!q_b_103),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~2 .extended_lut = "off";
defparam \ram_data_out2~2 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~2 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~2 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_104),
	.datad(!q_b_105),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~2 .extended_lut = "off";
defparam \ram_data_out3~2 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~2 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~2 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_106),
	.datad(!q_b_107),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~2 .extended_lut = "off";
defparam \ram_data_out0~2 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~2 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~3 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_11),
	.datad(!q_b_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~3 .extended_lut = "off";
defparam \ram_data_out1~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~3 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~3 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_112),
	.datad(!q_b_113),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~3 .extended_lut = "off";
defparam \ram_data_out2~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~3 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~3 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_114),
	.datad(!q_b_115),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~3 .extended_lut = "off";
defparam \ram_data_out3~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~3 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~3 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_116),
	.datad(!q_b_117),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~3 .extended_lut = "off";
defparam \ram_data_out0~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~3 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~4 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_12),
	.datad(!q_b_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~4 .extended_lut = "off";
defparam \ram_data_out1~4 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~4 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~4 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_122),
	.datad(!q_b_123),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~4 .extended_lut = "off";
defparam \ram_data_out2~4 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~4 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~4 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_124),
	.datad(!q_b_125),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~4 .extended_lut = "off";
defparam \ram_data_out3~4 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~4 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~4 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_126),
	.datad(!q_b_127),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~4 .extended_lut = "off";
defparam \ram_data_out0~4 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~4 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~5 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_15),
	.datad(!q_b_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~5 .extended_lut = "off";
defparam \ram_data_out1~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~5 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~5 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_152),
	.datad(!q_b_153),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~5 .extended_lut = "off";
defparam \ram_data_out2~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~5 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~5 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_154),
	.datad(!q_b_155),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~5 .extended_lut = "off";
defparam \ram_data_out3~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~5 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~5 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_156),
	.datad(!q_b_157),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~5 .extended_lut = "off";
defparam \ram_data_out0~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~5 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~6 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_7),
	.datad(!q_b_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~6 .extended_lut = "off";
defparam \ram_data_out1~6 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~6 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~6 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_72),
	.datad(!q_b_73),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~6 .extended_lut = "off";
defparam \ram_data_out2~6 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~6 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~6 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_74),
	.datad(!q_b_75),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~6 .extended_lut = "off";
defparam \ram_data_out3~6 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~6 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~6 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_76),
	.datad(!q_b_77),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~6 .extended_lut = "off";
defparam \ram_data_out0~6 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~6 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~7 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_6),
	.datad(!q_b_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~7 .extended_lut = "off";
defparam \ram_data_out1~7 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~7 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~7 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_62),
	.datad(!q_b_63),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~7 .extended_lut = "off";
defparam \ram_data_out2~7 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~7 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~7 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_64),
	.datad(!q_b_65),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~7 .extended_lut = "off";
defparam \ram_data_out3~7 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~7 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~7 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_66),
	.datad(!q_b_67),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~7 .extended_lut = "off";
defparam \ram_data_out0~7 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~7 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~8 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_3),
	.datad(!q_b_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~8 .extended_lut = "off";
defparam \ram_data_out1~8 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~8 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~8 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_32),
	.datad(!q_b_33),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~8 .extended_lut = "off";
defparam \ram_data_out2~8 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~8 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~8 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_34),
	.datad(!q_b_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~8 .extended_lut = "off";
defparam \ram_data_out3~8 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~8 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~8 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_36),
	.datad(!q_b_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~8 .extended_lut = "off";
defparam \ram_data_out0~8 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~8 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~9 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_4),
	.datad(!q_b_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~9 .extended_lut = "off";
defparam \ram_data_out1~9 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~9 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~9 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_42),
	.datad(!q_b_43),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~9 .extended_lut = "off";
defparam \ram_data_out2~9 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~9 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~9 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_44),
	.datad(!q_b_45),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~9 .extended_lut = "off";
defparam \ram_data_out3~9 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~9 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~9 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_46),
	.datad(!q_b_47),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~9 .extended_lut = "off";
defparam \ram_data_out0~9 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~9 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~10 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_5),
	.datad(!q_b_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~10 .extended_lut = "off";
defparam \ram_data_out1~10 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~10 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~10 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_52),
	.datad(!q_b_53),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~10 .extended_lut = "off";
defparam \ram_data_out2~10 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~10 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~10 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_54),
	.datad(!q_b_55),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~10 .extended_lut = "off";
defparam \ram_data_out3~10 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~10 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~10 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_56),
	.datad(!q_b_57),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~10 .extended_lut = "off";
defparam \ram_data_out0~10 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~10 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~11 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_2),
	.datad(!q_b_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~11 .extended_lut = "off";
defparam \ram_data_out1~11 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~11 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~11 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_22),
	.datad(!q_b_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~11 .extended_lut = "off";
defparam \ram_data_out2~11 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~11 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~11 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_24),
	.datad(!q_b_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~11 .extended_lut = "off";
defparam \ram_data_out3~11 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~11 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~11 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_26),
	.datad(!q_b_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~11 .extended_lut = "off";
defparam \ram_data_out0~11 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~11 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~12 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_8),
	.datad(!q_b_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~12 .extended_lut = "off";
defparam \ram_data_out2~12 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~12 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~12 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_82),
	.datad(!q_b_83),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~12 .extended_lut = "off";
defparam \ram_data_out3~12 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~12 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~12 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_84),
	.datad(!q_b_85),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~12 .extended_lut = "off";
defparam \ram_data_out0~12 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~12 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~12 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_86),
	.datad(!q_b_87),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~12 .extended_lut = "off";
defparam \ram_data_out1~12 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~12 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~13 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_9),
	.datad(!q_b_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~13 .extended_lut = "off";
defparam \ram_data_out2~13 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~13 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~13 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_92),
	.datad(!q_b_93),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~13 .extended_lut = "off";
defparam \ram_data_out3~13 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~13 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~13 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_94),
	.datad(!q_b_95),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~13 .extended_lut = "off";
defparam \ram_data_out0~13 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~13 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~13 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_96),
	.datad(!q_b_97),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~13 .extended_lut = "off";
defparam \ram_data_out1~13 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~13 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~14 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_0),
	.datad(!q_b_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~14 .extended_lut = "off";
defparam \ram_data_out3~14 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~14 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~14 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_02),
	.datad(!q_b_03),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~14 .extended_lut = "off";
defparam \ram_data_out0~14 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~14 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~14 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_04),
	.datad(!q_b_05),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~14 .extended_lut = "off";
defparam \ram_data_out1~14 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~14 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~14 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_06),
	.datad(!q_b_07),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~14 .extended_lut = "off";
defparam \ram_data_out2~14 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~14 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out3~15 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_1),
	.datad(!q_b_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out3~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out3~15 .extended_lut = "off";
defparam \ram_data_out3~15 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out3~15 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out0~15 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_17),
	.datad(!q_b_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out0~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out0~15 .extended_lut = "off";
defparam \ram_data_out0~15 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out0~15 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out1~15 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_19),
	.datad(!q_b_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out1~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out1~15 .extended_lut = "off";
defparam \ram_data_out1~15 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out1~15 .shared_arith = "off";

cyclonev_lcell_comb \ram_data_out2~15 (
	.dataa(!ram_a_not_b_vec_10),
	.datab(!data_rdy_vec_10),
	.datac(!q_b_118),
	.datad(!q_b_119),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_data_out2~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_data_out2~15 .extended_lut = "off";
defparam \ram_data_out2~15 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ram_data_out2~15 .shared_arith = "off";

endmodule

module IFFT_asj_fft_cxb_addr (
	global_clock_enable,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_2_1,
	ram_in_reg_3_3,
	ram_in_reg_3_0,
	rd_addr_d_0,
	rd_addr_d_1,
	sw_0,
	sw_1,
	ram_in_reg_3_01,
	ram_in_reg_2_11,
	ram_in_reg_3_31,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_2_1;
output 	ram_in_reg_3_3;
output 	ram_in_reg_3_0;
input 	rd_addr_d_0;
input 	rd_addr_d_1;
input 	sw_0;
input 	sw_1;
output 	ram_in_reg_3_01;
output 	ram_in_reg_2_11;
output 	ram_in_reg_3_31;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_in_reg[1][2]~0_combout ;
wire \ram_in_reg[3][3]~1_combout ;
wire \Mux0~0_combout ;


dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(rd_addr_d_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(rd_addr_d_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\ram_in_reg[1][2]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\ram_in_reg[3][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

cyclonev_lcell_comb \ram_in_reg[0][3]~_wirecell (
	.dataa(!ram_in_reg_3_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ram_in_reg_3_01),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_in_reg[0][3]~_wirecell .extended_lut = "off";
defparam \ram_in_reg[0][3]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ram_in_reg[0][3]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \ram_in_reg[1][2]~_wirecell (
	.dataa(!ram_in_reg_2_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ram_in_reg_2_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_in_reg[1][2]~_wirecell .extended_lut = "off";
defparam \ram_in_reg[1][2]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ram_in_reg[1][2]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \ram_in_reg[3][3]~_wirecell (
	.dataa(!ram_in_reg_3_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ram_in_reg_3_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_in_reg[3][3]~_wirecell .extended_lut = "off";
defparam \ram_in_reg[3][3]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ram_in_reg[3][3]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \ram_in_reg[1][2]~0 (
	.dataa(!sw_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_in_reg[1][2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_in_reg[1][2]~0 .extended_lut = "off";
defparam \ram_in_reg[1][2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ram_in_reg[1][2]~0 .shared_arith = "off";

cyclonev_lcell_comb \ram_in_reg[3][3]~1 (
	.dataa(!sw_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_in_reg[3][3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_in_reg[3][3]~1 .extended_lut = "off";
defparam \ram_in_reg[3][3]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ram_in_reg[3][3]~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!sw_0),
	.datab(!sw_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h6666666666666666;
defparam \Mux0~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_cxb_addr_1 (
	ram_block6a0,
	ram_block6a1,
	ram_block6a01,
	ram_block6a11,
	global_clock_enable,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_1_1,
	ram_in_reg_1_2,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_0_01,
	ram_in_reg_0_11,
	ram_in_reg_1_31,
	ram_in_reg_1_11,
	ram_in_reg_1_21,
	ram_in_reg_1_01,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_block6a0;
output 	ram_block6a1;
input 	ram_block6a01;
input 	ram_block6a11;
input 	global_clock_enable;
output 	ram_in_reg_0_1;
output 	ram_in_reg_1_3;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_2;
input 	ram_in_reg_2_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_0_01;
input 	ram_in_reg_0_11;
input 	ram_in_reg_1_31;
input 	ram_in_reg_1_11;
input 	ram_in_reg_1_21;
input 	ram_in_reg_1_01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \sw_0_arr_rtl_0|auto_generated|op_2~0_combout ;
wire \sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~1_sumout ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[0]~q ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~2 ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~5_sumout ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~q ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~6 ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~9_sumout ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[2]~q ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~10 ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~13_sumout ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[3]~q ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~14 ;
wire \sw_0_arr_rtl_0|auto_generated|op_1~17_sumout ;
wire \sw_0_arr_rtl_0|auto_generated|dffe3a[4]~q ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~1_sumout ;
wire \sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~2 ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~5_sumout ;
wire \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~q ;
wire \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~6 ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~9_sumout ;
wire \sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~10 ;
wire \sw_3_arr_rtl_0|auto_generated|op_1~13_sumout ;
wire \sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ;
wire \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout ;
wire \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout ;
wire \Mux7~0_combout ;
wire \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ;
wire \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ;
wire \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ;
wire \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ;
wire \Mux14~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;
wire \Mux6~0_combout ;
wire \Mux10~0_combout ;

wire [143:0] \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0_PORTBDATAOUT_bus ;
wire [143:0] \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1_PORTBDATAOUT_bus ;
wire [143:0] \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4_PORTBDATAOUT_bus ;
wire [143:0] \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2_PORTBDATAOUT_bus ;
wire [143:0] \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0_PORTBDATAOUT_bus ;
wire [143:0] \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3_PORTBDATAOUT_bus ;
wire [143:0] \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1_PORTBDATAOUT_bus ;
wire [143:0] \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5_PORTBDATAOUT_bus ;

assign ram_block6a0 = \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0_PORTBDATAOUT_bus [0];

assign ram_block6a1 = \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1_PORTBDATAOUT_bus [0];

assign \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout  = \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4_PORTBDATAOUT_bus [0];

assign \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout  = \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2_PORTBDATAOUT_bus [0];

assign \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout  = \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0_PORTBDATAOUT_bus [0];

assign \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout  = \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3_PORTBDATAOUT_bus [0];

assign \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout  = \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1_PORTBDATAOUT_bus [0];

assign \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout  = \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5_PORTBDATAOUT_bus [0];

cyclonev_ram_block \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_2_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,
\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|dffe3a[4]~q ,\sw_0_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_0_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,
\sw_0_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .clk1_output_clock_enable = "ena1";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_0|shift_taps_agv:auto_generated|altsyncram_pr91:altsyncram5|ALTSYNCRAM";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_address_width = 5;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_first_bit_number = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_last_address = 16;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_logical_ram_depth = 17;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_address_width = 5;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_data_out_clock = "clock1";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_first_bit_number = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_last_address = 16;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_logical_ram_depth = 17;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a0 .ram_block_type = "auto";

cyclonev_ram_block \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_3_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,
\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_0_arr_rtl_0|auto_generated|dffe3a[4]~q ,\sw_0_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_0_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,
\sw_0_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .clk0_core_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .clk0_input_clock_enable = "ena0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .clk1_output_clock_enable = "ena1";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .data_interleave_offset_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .data_interleave_width_in_bits = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_0_arr_rtl_0|shift_taps_agv:auto_generated|altsyncram_pr91:altsyncram5|ALTSYNCRAM";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .operation_mode = "dual_port";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_address_width = 5;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_data_out_clock = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_first_bit_number = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_last_address = 16;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_logical_ram_depth = 17;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_address_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_address_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_address_width = 5;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_data_out_clear = "none";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_data_out_clock = "clock1";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_data_width = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_first_address = 0;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_first_bit_number = 1;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_last_address = 16;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_logical_ram_depth = 17;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_logical_ram_width = 2;
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_read_enable_clock = "clock0";
defparam \sw_0_arr_rtl_0|auto_generated|altsyncram5|ram_block6a1 .ram_block_type = "auto";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .lut_mask = 64'h0000000000000000;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .shared_arith = "off";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sw_0_arr_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|op_2~0 (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|op_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|op_2~0 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|op_2~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \sw_0_arr_rtl_0|auto_generated|op_2~0 .shared_arith = "off";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0 (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0 .lut_mask = 64'hFFFFBFFFFFFFBFFF;
defparam \sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0 .shared_arith = "off";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|op_1~1 (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(!\sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h000055FF000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|dffe3a[0] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|dffe3a[1] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|dffe3a[2] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(\sw_0_arr_rtl_0|auto_generated|op_1~14 ),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|dffe3a[3] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_lcell_comb \sw_0_arr_rtl_0|auto_generated|op_1~17 (
	.dataa(!\sw_0_arr_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_0_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(!\sw_0_arr_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\sw_0_arr_rtl_0|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_0_arr_rtl_0|auto_generated|op_1~17_sumout ),
	.cout(),
	.shareout());
defparam \sw_0_arr_rtl_0|auto_generated|op_1~17 .extended_lut = "off";
defparam \sw_0_arr_rtl_0|auto_generated|op_1~17 .lut_mask = 64'h0000FFAA000000FF;
defparam \sw_0_arr_rtl_0|auto_generated|op_1~17 .shared_arith = "off";

dffeas \sw_0_arr_rtl_0|auto_generated|dffe3a[4] (
	.clk(clk),
	.d(\sw_0_arr_rtl_0|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_0_arr_rtl_0|auto_generated|dffe3a[4]~q ),
	.prn(vcc));
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \sw_0_arr_rtl_0|auto_generated|dffe3a[4] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\sw_3_arr_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|dffe3a[0] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_3_arr_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\sw_3_arr_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\sw_3_arr_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|dffe3a[1] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_3_arr_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\sw_3_arr_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|dffe3a[2] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \sw_3_arr_rtl_0|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\sw_3_arr_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\sw_3_arr_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(),
	.shareout());
defparam \sw_3_arr_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \sw_3_arr_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \sw_3_arr_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \sw_3_arr_rtl_0|auto_generated|dffe3a[3] (
	.clk(clk),
	.d(\sw_3_arr_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \sw_3_arr_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_ram_block \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_0_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .clk0_core_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .clk0_input_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .clk1_output_clock_enable = "ena1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .data_interleave_offset_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .data_interleave_width_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_3_arr_rtl_0|shift_taps_egv:auto_generated|altsyncram_tr91:altsyncram4|ALTSYNCRAM";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .operation_mode = "dual_port";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_data_out_clock = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_first_bit_number = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_address_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_data_out_clock = "clock1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_first_bit_number = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_read_enable_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4 .ram_block_type = "auto";

cyclonev_ram_block \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_0_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .clk0_core_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .clk0_input_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .clk1_output_clock_enable = "ena1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .data_interleave_offset_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .data_interleave_width_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_3_arr_rtl_0|shift_taps_egv:auto_generated|altsyncram_tr91:altsyncram4|ALTSYNCRAM";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .operation_mode = "dual_port";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_data_out_clock = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_first_bit_number = 2;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_address_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_data_out_clock = "clock1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_first_bit_number = 2;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_read_enable_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2 .ram_block_type = "auto";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!ram_block6a01),
	.datab(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout ),
	.datac(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h2727272727272727;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_ram_block \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_31}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .clk0_core_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .clk0_input_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .clk1_output_clock_enable = "ena1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .data_interleave_offset_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .data_interleave_width_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_3_arr_rtl_0|shift_taps_egv:auto_generated|altsyncram_tr91:altsyncram4|ALTSYNCRAM";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .operation_mode = "dual_port";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_data_out_clock = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_first_bit_number = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_address_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_data_out_clock = "clock1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_first_bit_number = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_read_enable_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0 .ram_block_type = "auto";

cyclonev_ram_block \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .clk0_core_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .clk0_input_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .clk1_output_clock_enable = "ena1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .data_interleave_offset_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .data_interleave_width_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_3_arr_rtl_0|shift_taps_egv:auto_generated|altsyncram_tr91:altsyncram4|ALTSYNCRAM";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .operation_mode = "dual_port";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_data_out_clock = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_first_bit_number = 3;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_address_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_data_out_clock = "clock1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_first_bit_number = 3;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_read_enable_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3 .ram_block_type = "auto";

cyclonev_ram_block \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_21}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .clk0_core_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .clk0_input_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .clk1_output_clock_enable = "ena1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .data_interleave_offset_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .data_interleave_width_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_3_arr_rtl_0|shift_taps_egv:auto_generated|altsyncram_tr91:altsyncram4|ALTSYNCRAM";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .operation_mode = "dual_port";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_data_out_clock = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_first_bit_number = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_address_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_data_out_clock = "clock1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_first_bit_number = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_read_enable_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1 .ram_block_type = "auto";

cyclonev_ram_block \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ram_in_reg_1_01}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\sw_3_arr_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\sw_3_arr_rtl_0|auto_generated|dffe3a[3]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[2]~q ,\sw_3_arr_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\sw_3_arr_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .clk0_core_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .clk0_input_clock_enable = "ena0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .clk1_output_clock_enable = "ena1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .data_interleave_offset_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .data_interleave_width_in_bits = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_cxb_addr:\\gen_wrsw_1:ram_cxb_wr|altshift_taps:sw_3_arr_rtl_0|shift_taps_egv:auto_generated|altsyncram_tr91:altsyncram4|ALTSYNCRAM";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .mixed_port_feed_through_mode = "dont_care";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .operation_mode = "dual_port";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_data_out_clock = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_first_bit_number = 5;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_address_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_address_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_address_width = 4;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_data_out_clear = "none";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_data_out_clock = "clock1";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_data_width = 1;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_first_address = 0;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_first_bit_number = 5;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_last_address = 15;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_logical_ram_depth = 16;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_logical_ram_width = 6;
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_read_enable_clock = "clock0";
defparam \sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5 .ram_block_type = "auto";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ),
	.datab(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ),
	.datac(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ),
	.datad(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ),
	.datae(!ram_block6a11),
	.dataf(!ram_block6a01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!ram_block6a01),
	.datab(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout ),
	.datac(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h2727272727272727;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ),
	.datab(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ),
	.datac(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ),
	.datad(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ),
	.datae(!ram_block6a11),
	.dataf(!ram_block6a01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ),
	.datab(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ),
	.datac(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ),
	.datad(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ),
	.datae(!ram_block6a11),
	.dataf(!ram_block6a01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ),
	.datab(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ),
	.datac(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ),
	.datad(!\sw_3_arr_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ),
	.datae(!ram_block6a11),
	.dataf(!ram_block6a01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_cxb_addr_2 (
	global_clock_enable,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_0_0,
	ram_in_reg_0_1,
	ram_in_reg_1_3,
	ram_in_reg_1_1,
	ram_in_reg_1_2,
	ram_in_reg_1_0,
	rd_addr_d_2,
	rd_addr_d_3,
	rd_addr_d_0,
	sw_0,
	rd_addr_c_0,
	rd_addr_b_1,
	sw_1,
	rd_addr_d_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_0_0;
output 	ram_in_reg_0_1;
output 	ram_in_reg_1_3;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_0;
input 	rd_addr_d_2;
input 	rd_addr_d_3;
input 	rd_addr_d_0;
input 	sw_0;
input 	rd_addr_c_0;
input 	rd_addr_b_1;
input 	sw_1;
input 	rd_addr_d_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux3~0_combout ;
wire \Mux7~0_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux10~0_combout ;
wire \Mux2~0_combout ;


dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(rd_addr_d_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(rd_addr_d_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux14~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!rd_addr_d_0),
	.datab(!sw_0),
	.datac(!rd_addr_c_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h4747474747474747;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!rd_addr_d_0),
	.datab(!sw_0),
	.datac(!rd_addr_c_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h4747474747474747;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!rd_addr_b_1),
	.datab(!sw_1),
	.datac(!rd_addr_d_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h4747474747474747;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~1 (
	.dataa(!rd_addr_b_1),
	.datab(!sw_1),
	.datac(!rd_addr_d_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~1 .extended_lut = "off";
defparam \Mux14~1 .lut_mask = 64'h4747474747474747;
defparam \Mux14~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!sw_0),
	.datab(!\Mux14~0_combout ),
	.datac(!\Mux14~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h2727272727272727;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!sw_0),
	.datab(!\Mux14~0_combout ),
	.datac(!\Mux14~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h2727272727272727;
defparam \Mux2~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_cxb_data (
	reg_no_twiddle603,
	reg_no_twiddle607,
	reg_no_twiddle617,
	reg_no_twiddle613,
	reg_no_twiddle604,
	reg_no_twiddle614,
	reg_no_twiddle605,
	reg_no_twiddle615,
	reg_no_twiddle606,
	reg_no_twiddle616,
	reg_no_twiddle602,
	ram_block6a3,
	ram_block6a2,
	reg_no_twiddle612,
	reg_no_twiddle601,
	reg_no_twiddle611,
	reg_no_twiddle600,
	reg_no_twiddle610,
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_3_11,
	tdl_arr_7_11,
	tdl_arr_3_12,
	tdl_arr_7_12,
	tdl_arr_3_13,
	tdl_arr_7_13,
	tdl_arr_3_14,
	tdl_arr_7_14,
	tdl_arr_3_15,
	tdl_arr_7_15,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_4_12,
	tdl_arr_4_13,
	tdl_arr_4_14,
	tdl_arr_4_15,
	tdl_arr_5_1,
	tdl_arr_5_11,
	tdl_arr_5_12,
	tdl_arr_5_13,
	tdl_arr_5_14,
	tdl_arr_5_15,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_6_12,
	tdl_arr_6_13,
	tdl_arr_6_14,
	tdl_arr_6_15,
	ram_in_reg_2_3,
	ram_in_reg_2_0,
	ram_in_reg_2_1,
	ram_in_reg_2_2,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_5,
	ram_in_reg_2_6,
	ram_in_reg_3_3,
	ram_in_reg_3_0,
	ram_in_reg_3_1,
	ram_in_reg_3_2,
	ram_in_reg_3_7,
	ram_in_reg_3_4,
	ram_in_reg_3_5,
	ram_in_reg_3_6,
	ram_in_reg_4_3,
	ram_in_reg_4_0,
	ram_in_reg_4_1,
	ram_in_reg_4_2,
	ram_in_reg_4_7,
	ram_in_reg_4_4,
	ram_in_reg_4_5,
	ram_in_reg_4_6,
	ram_in_reg_5_3,
	ram_in_reg_5_0,
	ram_in_reg_5_1,
	ram_in_reg_5_2,
	ram_in_reg_5_7,
	ram_in_reg_5_4,
	ram_in_reg_5_5,
	ram_in_reg_5_6,
	ram_in_reg_6_3,
	ram_in_reg_6_0,
	ram_in_reg_6_1,
	ram_in_reg_6_2,
	ram_in_reg_6_7,
	ram_in_reg_6_4,
	ram_in_reg_6_5,
	ram_in_reg_6_6,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_1,
	ram_in_reg_7_2,
	ram_in_reg_7_7,
	ram_in_reg_7_4,
	ram_in_reg_7_5,
	ram_in_reg_7_6,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_2_12,
	tdl_arr_2_13,
	tdl_arr_2_14,
	tdl_arr_2_15,
	ram_in_reg_1_3,
	ram_in_reg_1_0,
	ram_in_reg_1_1,
	ram_in_reg_1_2,
	ram_in_reg_1_7,
	ram_in_reg_1_4,
	ram_in_reg_1_5,
	ram_in_reg_1_6,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_1_12,
	tdl_arr_1_13,
	tdl_arr_1_14,
	tdl_arr_1_15,
	ram_in_reg_0_3,
	ram_in_reg_0_0,
	ram_in_reg_0_1,
	ram_in_reg_0_2,
	ram_in_reg_0_7,
	ram_in_reg_0_4,
	ram_in_reg_0_5,
	ram_in_reg_0_6,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_0_12,
	tdl_arr_0_13,
	tdl_arr_0_14,
	tdl_arr_0_15,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reg_no_twiddle603;
input 	reg_no_twiddle607;
input 	reg_no_twiddle617;
input 	reg_no_twiddle613;
input 	reg_no_twiddle604;
input 	reg_no_twiddle614;
input 	reg_no_twiddle605;
input 	reg_no_twiddle615;
input 	reg_no_twiddle606;
input 	reg_no_twiddle616;
input 	reg_no_twiddle602;
input 	ram_block6a3;
input 	ram_block6a2;
input 	reg_no_twiddle612;
input 	reg_no_twiddle601;
input 	reg_no_twiddle611;
input 	reg_no_twiddle600;
input 	reg_no_twiddle610;
input 	global_clock_enable;
input 	tdl_arr_3_1;
input 	tdl_arr_7_1;
input 	tdl_arr_3_11;
input 	tdl_arr_7_11;
input 	tdl_arr_3_12;
input 	tdl_arr_7_12;
input 	tdl_arr_3_13;
input 	tdl_arr_7_13;
input 	tdl_arr_3_14;
input 	tdl_arr_7_14;
input 	tdl_arr_3_15;
input 	tdl_arr_7_15;
input 	tdl_arr_4_1;
input 	tdl_arr_4_11;
input 	tdl_arr_4_12;
input 	tdl_arr_4_13;
input 	tdl_arr_4_14;
input 	tdl_arr_4_15;
input 	tdl_arr_5_1;
input 	tdl_arr_5_11;
input 	tdl_arr_5_12;
input 	tdl_arr_5_13;
input 	tdl_arr_5_14;
input 	tdl_arr_5_15;
input 	tdl_arr_6_1;
input 	tdl_arr_6_11;
input 	tdl_arr_6_12;
input 	tdl_arr_6_13;
input 	tdl_arr_6_14;
input 	tdl_arr_6_15;
output 	ram_in_reg_2_3;
output 	ram_in_reg_2_0;
output 	ram_in_reg_2_1;
output 	ram_in_reg_2_2;
output 	ram_in_reg_2_7;
output 	ram_in_reg_2_4;
output 	ram_in_reg_2_5;
output 	ram_in_reg_2_6;
output 	ram_in_reg_3_3;
output 	ram_in_reg_3_0;
output 	ram_in_reg_3_1;
output 	ram_in_reg_3_2;
output 	ram_in_reg_3_7;
output 	ram_in_reg_3_4;
output 	ram_in_reg_3_5;
output 	ram_in_reg_3_6;
output 	ram_in_reg_4_3;
output 	ram_in_reg_4_0;
output 	ram_in_reg_4_1;
output 	ram_in_reg_4_2;
output 	ram_in_reg_4_7;
output 	ram_in_reg_4_4;
output 	ram_in_reg_4_5;
output 	ram_in_reg_4_6;
output 	ram_in_reg_5_3;
output 	ram_in_reg_5_0;
output 	ram_in_reg_5_1;
output 	ram_in_reg_5_2;
output 	ram_in_reg_5_7;
output 	ram_in_reg_5_4;
output 	ram_in_reg_5_5;
output 	ram_in_reg_5_6;
output 	ram_in_reg_6_3;
output 	ram_in_reg_6_0;
output 	ram_in_reg_6_1;
output 	ram_in_reg_6_2;
output 	ram_in_reg_6_7;
output 	ram_in_reg_6_4;
output 	ram_in_reg_6_5;
output 	ram_in_reg_6_6;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_0;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_7;
output 	ram_in_reg_7_4;
output 	ram_in_reg_7_5;
output 	ram_in_reg_7_6;
input 	tdl_arr_2_1;
input 	tdl_arr_2_11;
input 	tdl_arr_2_12;
input 	tdl_arr_2_13;
input 	tdl_arr_2_14;
input 	tdl_arr_2_15;
output 	ram_in_reg_1_3;
output 	ram_in_reg_1_0;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_7;
output 	ram_in_reg_1_4;
output 	ram_in_reg_1_5;
output 	ram_in_reg_1_6;
input 	tdl_arr_1_1;
input 	tdl_arr_1_11;
input 	tdl_arr_1_12;
input 	tdl_arr_1_13;
input 	tdl_arr_1_14;
input 	tdl_arr_1_15;
output 	ram_in_reg_0_3;
output 	ram_in_reg_0_0;
output 	ram_in_reg_0_1;
output 	ram_in_reg_0_2;
output 	ram_in_reg_0_7;
output 	ram_in_reg_0_4;
output 	ram_in_reg_0_5;
output 	ram_in_reg_0_6;
input 	tdl_arr_0_1;
input 	tdl_arr_0_11;
input 	tdl_arr_0_12;
input 	tdl_arr_0_13;
input 	tdl_arr_0_14;
input 	tdl_arr_0_15;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux29~0_combout ;
wire \Mux5~0_combout ;
wire \Mux13~0_combout ;
wire \Mux21~0_combout ;
wire \Mux61~0_combout ;
wire \Mux37~0_combout ;
wire \Mux45~0_combout ;
wire \Mux53~0_combout ;
wire \Mux28~0_combout ;
wire \Mux4~0_combout ;
wire \Mux12~0_combout ;
wire \Mux20~0_combout ;
wire \Mux60~0_combout ;
wire \Mux36~0_combout ;
wire \Mux44~0_combout ;
wire \Mux52~0_combout ;
wire \Mux27~0_combout ;
wire \Mux3~0_combout ;
wire \Mux11~0_combout ;
wire \Mux19~0_combout ;
wire \Mux59~0_combout ;
wire \Mux35~0_combout ;
wire \Mux43~0_combout ;
wire \Mux51~0_combout ;
wire \Mux26~0_combout ;
wire \Mux2~0_combout ;
wire \Mux10~0_combout ;
wire \Mux18~0_combout ;
wire \Mux58~0_combout ;
wire \Mux34~0_combout ;
wire \Mux42~0_combout ;
wire \Mux50~0_combout ;
wire \Mux25~0_combout ;
wire \Mux1~0_combout ;
wire \Mux9~0_combout ;
wire \Mux17~0_combout ;
wire \Mux57~0_combout ;
wire \Mux33~0_combout ;
wire \Mux41~0_combout ;
wire \Mux49~0_combout ;
wire \Mux24~0_combout ;
wire \Mux0~0_combout ;
wire \Mux8~0_combout ;
wire \Mux16~0_combout ;
wire \Mux56~0_combout ;
wire \Mux32~0_combout ;
wire \Mux40~0_combout ;
wire \Mux48~0_combout ;
wire \Mux30~0_combout ;
wire \Mux6~0_combout ;
wire \Mux14~0_combout ;
wire \Mux22~0_combout ;
wire \Mux62~0_combout ;
wire \Mux38~0_combout ;
wire \Mux46~0_combout ;
wire \Mux54~0_combout ;
wire \Mux31~0_combout ;
wire \Mux7~0_combout ;
wire \Mux15~0_combout ;
wire \Mux23~0_combout ;
wire \Mux63~0_combout ;
wire \Mux39~0_combout ;
wire \Mux47~0_combout ;
wire \Mux55~0_combout ;


dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\Mux29~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\Mux21~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\Mux61~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\Mux45~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\Mux53~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\Mux28~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\Mux20~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\Mux60~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\Mux36~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\Mux44~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\Mux52~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\Mux27~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\Mux19~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\Mux59~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\Mux35~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\Mux43~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\Mux51~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\Mux26~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\Mux18~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\Mux58~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\Mux34~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\Mux42~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\Mux50~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\Mux25~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\Mux57~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\Mux33~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\Mux41~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\Mux49~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\Mux24~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\Mux16~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\Mux56~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\Mux32~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\Mux40~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\Mux48~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux30~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux22~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\Mux62~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\Mux38~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\Mux46~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\Mux54~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\Mux31~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\Mux23~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\Mux63~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\Mux39~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\Mux47~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\Mux55~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

cyclonev_lcell_comb \Mux29~0 (
	.dataa(!tdl_arr_2_1),
	.datab(!tdl_arr_2_11),
	.datac(!tdl_arr_2_12),
	.datad(!reg_no_twiddle602),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux29~0 .extended_lut = "off";
defparam \Mux29~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux29~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!reg_no_twiddle602),
	.datab(!tdl_arr_2_12),
	.datac(!tdl_arr_2_1),
	.datad(!tdl_arr_2_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux5~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!tdl_arr_2_11),
	.datab(!tdl_arr_2_1),
	.datac(!reg_no_twiddle602),
	.datad(!tdl_arr_2_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "off";
defparam \Mux13~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux13~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux21~0 (
	.dataa(!tdl_arr_2_12),
	.datab(!reg_no_twiddle602),
	.datac(!tdl_arr_2_11),
	.datad(!tdl_arr_2_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux21~0 .extended_lut = "off";
defparam \Mux21~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux21~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux61~0 (
	.dataa(!tdl_arr_2_13),
	.datab(!tdl_arr_2_14),
	.datac(!tdl_arr_2_15),
	.datad(!reg_no_twiddle612),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux61~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux61~0 .extended_lut = "off";
defparam \Mux61~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux61~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!reg_no_twiddle612),
	.datab(!tdl_arr_2_15),
	.datac(!tdl_arr_2_13),
	.datad(!tdl_arr_2_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux37~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~0 (
	.dataa(!tdl_arr_2_14),
	.datab(!tdl_arr_2_13),
	.datac(!reg_no_twiddle612),
	.datad(!tdl_arr_2_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~0 .extended_lut = "off";
defparam \Mux45~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux53~0 (
	.dataa(!tdl_arr_2_15),
	.datab(!reg_no_twiddle612),
	.datac(!tdl_arr_2_14),
	.datad(!tdl_arr_2_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux53~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux53~0 .extended_lut = "off";
defparam \Mux53~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux53~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux28~0 (
	.dataa(!tdl_arr_3_14),
	.datab(!tdl_arr_3_13),
	.datac(!tdl_arr_3_11),
	.datad(!reg_no_twiddle603),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux28~0 .extended_lut = "off";
defparam \Mux28~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux28~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!reg_no_twiddle603),
	.datab(!tdl_arr_3_11),
	.datac(!tdl_arr_3_14),
	.datad(!tdl_arr_3_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!tdl_arr_3_13),
	.datab(!tdl_arr_3_14),
	.datac(!reg_no_twiddle603),
	.datad(!tdl_arr_3_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "off";
defparam \Mux12~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux12~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux20~0 (
	.dataa(!tdl_arr_3_11),
	.datab(!reg_no_twiddle603),
	.datac(!tdl_arr_3_13),
	.datad(!tdl_arr_3_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux20~0 .extended_lut = "off";
defparam \Mux20~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux20~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux60~0 (
	.dataa(!tdl_arr_3_15),
	.datab(!tdl_arr_3_1),
	.datac(!tdl_arr_3_12),
	.datad(!reg_no_twiddle613),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux60~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux60~0 .extended_lut = "off";
defparam \Mux60~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux60~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux36~0 (
	.dataa(!reg_no_twiddle613),
	.datab(!tdl_arr_3_12),
	.datac(!tdl_arr_3_15),
	.datad(!tdl_arr_3_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux36~0 .extended_lut = "off";
defparam \Mux36~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux36~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~0 (
	.dataa(!tdl_arr_3_1),
	.datab(!tdl_arr_3_15),
	.datac(!reg_no_twiddle613),
	.datad(!tdl_arr_3_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~0 .extended_lut = "off";
defparam \Mux44~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux52~0 (
	.dataa(!tdl_arr_3_12),
	.datab(!reg_no_twiddle613),
	.datac(!tdl_arr_3_1),
	.datad(!tdl_arr_3_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux52~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux52~0 .extended_lut = "off";
defparam \Mux52~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux52~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!tdl_arr_4_14),
	.datab(!tdl_arr_4_13),
	.datac(!tdl_arr_4_11),
	.datad(!reg_no_twiddle604),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!reg_no_twiddle604),
	.datab(!tdl_arr_4_11),
	.datac(!tdl_arr_4_14),
	.datad(!tdl_arr_4_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!tdl_arr_4_13),
	.datab(!tdl_arr_4_14),
	.datac(!reg_no_twiddle604),
	.datad(!tdl_arr_4_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!tdl_arr_4_11),
	.datab(!reg_no_twiddle604),
	.datac(!tdl_arr_4_13),
	.datad(!tdl_arr_4_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux59~0 (
	.dataa(!tdl_arr_4_15),
	.datab(!tdl_arr_4_1),
	.datac(!tdl_arr_4_12),
	.datad(!reg_no_twiddle614),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux59~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux59~0 .extended_lut = "off";
defparam \Mux59~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux59~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~0 (
	.dataa(!reg_no_twiddle614),
	.datab(!tdl_arr_4_12),
	.datac(!tdl_arr_4_15),
	.datad(!tdl_arr_4_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~0 .extended_lut = "off";
defparam \Mux35~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux35~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~0 (
	.dataa(!tdl_arr_4_1),
	.datab(!tdl_arr_4_15),
	.datac(!reg_no_twiddle614),
	.datad(!tdl_arr_4_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~0 .extended_lut = "off";
defparam \Mux43~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux51~0 (
	.dataa(!tdl_arr_4_12),
	.datab(!reg_no_twiddle614),
	.datac(!tdl_arr_4_1),
	.datad(!tdl_arr_4_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux51~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux51~0 .extended_lut = "off";
defparam \Mux51~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux51~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!tdl_arr_5_14),
	.datab(!tdl_arr_5_13),
	.datac(!tdl_arr_5_11),
	.datad(!reg_no_twiddle605),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!reg_no_twiddle605),
	.datab(!tdl_arr_5_11),
	.datac(!tdl_arr_5_14),
	.datad(!tdl_arr_5_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!tdl_arr_5_13),
	.datab(!tdl_arr_5_14),
	.datac(!reg_no_twiddle605),
	.datad(!tdl_arr_5_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!tdl_arr_5_11),
	.datab(!reg_no_twiddle605),
	.datac(!tdl_arr_5_13),
	.datad(!tdl_arr_5_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "off";
defparam \Mux18~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux58~0 (
	.dataa(!tdl_arr_5_15),
	.datab(!tdl_arr_5_1),
	.datac(!tdl_arr_5_12),
	.datad(!reg_no_twiddle615),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux58~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux58~0 .extended_lut = "off";
defparam \Mux58~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux58~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~0 (
	.dataa(!reg_no_twiddle615),
	.datab(!tdl_arr_5_12),
	.datac(!tdl_arr_5_15),
	.datad(!tdl_arr_5_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~0 .extended_lut = "off";
defparam \Mux34~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux34~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~0 (
	.dataa(!tdl_arr_5_1),
	.datab(!tdl_arr_5_15),
	.datac(!reg_no_twiddle615),
	.datad(!tdl_arr_5_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~0 .extended_lut = "off";
defparam \Mux42~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux50~0 (
	.dataa(!tdl_arr_5_12),
	.datab(!reg_no_twiddle615),
	.datac(!tdl_arr_5_1),
	.datad(!tdl_arr_5_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux50~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux50~0 .extended_lut = "off";
defparam \Mux50~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux50~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!tdl_arr_6_14),
	.datab(!tdl_arr_6_13),
	.datac(!tdl_arr_6_11),
	.datad(!reg_no_twiddle606),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!reg_no_twiddle606),
	.datab(!tdl_arr_6_11),
	.datac(!tdl_arr_6_14),
	.datad(!tdl_arr_6_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!tdl_arr_6_13),
	.datab(!tdl_arr_6_14),
	.datac(!reg_no_twiddle606),
	.datad(!tdl_arr_6_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!tdl_arr_6_11),
	.datab(!reg_no_twiddle606),
	.datac(!tdl_arr_6_13),
	.datad(!tdl_arr_6_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "off";
defparam \Mux17~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux57~0 (
	.dataa(!tdl_arr_6_15),
	.datab(!tdl_arr_6_1),
	.datac(!tdl_arr_6_12),
	.datad(!reg_no_twiddle616),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux57~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux57~0 .extended_lut = "off";
defparam \Mux57~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux57~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~0 (
	.dataa(!reg_no_twiddle616),
	.datab(!tdl_arr_6_12),
	.datac(!tdl_arr_6_15),
	.datad(!tdl_arr_6_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~0 .extended_lut = "off";
defparam \Mux33~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux33~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~0 (
	.dataa(!tdl_arr_6_1),
	.datab(!tdl_arr_6_15),
	.datac(!reg_no_twiddle616),
	.datad(!tdl_arr_6_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~0 .extended_lut = "off";
defparam \Mux41~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux49~0 (
	.dataa(!tdl_arr_6_12),
	.datab(!reg_no_twiddle616),
	.datac(!tdl_arr_6_1),
	.datad(!tdl_arr_6_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux49~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux49~0 .extended_lut = "off";
defparam \Mux49~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux49~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!tdl_arr_7_14),
	.datab(!tdl_arr_7_13),
	.datac(!tdl_arr_7_11),
	.datad(!reg_no_twiddle607),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!reg_no_twiddle607),
	.datab(!tdl_arr_7_11),
	.datac(!tdl_arr_7_14),
	.datad(!tdl_arr_7_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!tdl_arr_7_13),
	.datab(!tdl_arr_7_14),
	.datac(!reg_no_twiddle607),
	.datad(!tdl_arr_7_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!tdl_arr_7_11),
	.datab(!reg_no_twiddle607),
	.datac(!tdl_arr_7_13),
	.datad(!tdl_arr_7_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "off";
defparam \Mux16~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux16~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~0 (
	.dataa(!tdl_arr_7_15),
	.datab(!tdl_arr_7_1),
	.datac(!tdl_arr_7_12),
	.datad(!reg_no_twiddle617),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~0 .extended_lut = "off";
defparam \Mux56~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux56~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~0 (
	.dataa(!reg_no_twiddle617),
	.datab(!tdl_arr_7_12),
	.datac(!tdl_arr_7_15),
	.datad(!tdl_arr_7_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~0 .extended_lut = "off";
defparam \Mux32~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux32~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~0 (
	.dataa(!tdl_arr_7_1),
	.datab(!tdl_arr_7_15),
	.datac(!reg_no_twiddle617),
	.datad(!tdl_arr_7_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~0 .extended_lut = "off";
defparam \Mux40~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~0 (
	.dataa(!tdl_arr_7_12),
	.datab(!reg_no_twiddle617),
	.datac(!tdl_arr_7_1),
	.datad(!tdl_arr_7_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~0 .extended_lut = "off";
defparam \Mux48~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux48~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux30~0 (
	.dataa(!tdl_arr_1_1),
	.datab(!tdl_arr_1_11),
	.datac(!tdl_arr_1_12),
	.datad(!reg_no_twiddle601),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux30~0 .extended_lut = "off";
defparam \Mux30~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux30~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!reg_no_twiddle601),
	.datab(!tdl_arr_1_12),
	.datac(!tdl_arr_1_1),
	.datad(!tdl_arr_1_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!tdl_arr_1_11),
	.datab(!tdl_arr_1_1),
	.datac(!reg_no_twiddle601),
	.datad(!tdl_arr_1_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux22~0 (
	.dataa(!tdl_arr_1_12),
	.datab(!reg_no_twiddle601),
	.datac(!tdl_arr_1_11),
	.datad(!tdl_arr_1_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux22~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux62~0 (
	.dataa(!tdl_arr_1_13),
	.datab(!tdl_arr_1_14),
	.datac(!tdl_arr_1_15),
	.datad(!reg_no_twiddle611),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux62~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux62~0 .extended_lut = "off";
defparam \Mux62~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux62~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux38~0 (
	.dataa(!reg_no_twiddle611),
	.datab(!tdl_arr_1_15),
	.datac(!tdl_arr_1_13),
	.datad(!tdl_arr_1_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux38~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux38~0 .extended_lut = "off";
defparam \Mux38~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux38~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~0 (
	.dataa(!tdl_arr_1_14),
	.datab(!tdl_arr_1_13),
	.datac(!reg_no_twiddle611),
	.datad(!tdl_arr_1_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~0 .extended_lut = "off";
defparam \Mux46~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux54~0 (
	.dataa(!tdl_arr_1_15),
	.datab(!reg_no_twiddle611),
	.datac(!tdl_arr_1_14),
	.datad(!tdl_arr_1_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux54~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux54~0 .extended_lut = "off";
defparam \Mux54~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux54~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux31~0 (
	.dataa(!tdl_arr_0_1),
	.datab(!tdl_arr_0_11),
	.datac(!tdl_arr_0_12),
	.datad(!reg_no_twiddle600),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux31~0 .extended_lut = "off";
defparam \Mux31~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux31~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!reg_no_twiddle600),
	.datab(!tdl_arr_0_12),
	.datac(!tdl_arr_0_1),
	.datad(!tdl_arr_0_11),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!tdl_arr_0_11),
	.datab(!tdl_arr_0_1),
	.datac(!reg_no_twiddle600),
	.datad(!tdl_arr_0_12),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "off";
defparam \Mux15~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux15~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux23~0 (
	.dataa(!tdl_arr_0_12),
	.datab(!reg_no_twiddle600),
	.datac(!tdl_arr_0_11),
	.datad(!tdl_arr_0_1),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux23~0 .extended_lut = "off";
defparam \Mux23~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux23~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux63~0 (
	.dataa(!tdl_arr_0_13),
	.datab(!tdl_arr_0_14),
	.datac(!tdl_arr_0_15),
	.datad(!reg_no_twiddle610),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux63~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux63~0 .extended_lut = "off";
defparam \Mux63~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux63~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux39~0 (
	.dataa(!reg_no_twiddle610),
	.datab(!tdl_arr_0_15),
	.datac(!tdl_arr_0_13),
	.datad(!tdl_arr_0_14),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux39~0 .extended_lut = "off";
defparam \Mux39~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux39~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~0 (
	.dataa(!tdl_arr_0_14),
	.datab(!tdl_arr_0_13),
	.datac(!reg_no_twiddle610),
	.datad(!tdl_arr_0_15),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~0 .extended_lut = "off";
defparam \Mux47~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux55~0 (
	.dataa(!tdl_arr_0_15),
	.datab(!reg_no_twiddle610),
	.datac(!tdl_arr_0_14),
	.datad(!tdl_arr_0_13),
	.datae(!ram_block6a3),
	.dataf(!ram_block6a2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux55~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux55~0 .extended_lut = "off";
defparam \Mux55~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux55~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_cxb_data_r (
	lpp_ram_data_out_10_3,
	lpp_ram_data_out_10_0,
	lpp_ram_data_out_10_1,
	lpp_ram_data_out_10_2,
	tdl_arr_0_4,
	tdl_arr_1_4,
	lpp_ram_data_out_2_3,
	lpp_ram_data_out_2_0,
	lpp_ram_data_out_2_1,
	lpp_ram_data_out_2_2,
	lpp_ram_data_out_11_3,
	lpp_ram_data_out_11_0,
	lpp_ram_data_out_11_1,
	lpp_ram_data_out_11_2,
	lpp_ram_data_out_3_3,
	lpp_ram_data_out_3_0,
	lpp_ram_data_out_3_1,
	lpp_ram_data_out_3_2,
	lpp_ram_data_out_12_3,
	lpp_ram_data_out_12_0,
	lpp_ram_data_out_12_1,
	lpp_ram_data_out_12_2,
	lpp_ram_data_out_4_3,
	lpp_ram_data_out_4_0,
	lpp_ram_data_out_4_1,
	lpp_ram_data_out_4_2,
	lpp_ram_data_out_13_3,
	lpp_ram_data_out_13_0,
	lpp_ram_data_out_13_1,
	lpp_ram_data_out_13_2,
	lpp_ram_data_out_5_3,
	lpp_ram_data_out_5_0,
	lpp_ram_data_out_5_1,
	lpp_ram_data_out_5_2,
	lpp_ram_data_out_14_3,
	lpp_ram_data_out_14_0,
	lpp_ram_data_out_14_1,
	lpp_ram_data_out_14_2,
	lpp_ram_data_out_6_3,
	lpp_ram_data_out_6_0,
	lpp_ram_data_out_6_1,
	lpp_ram_data_out_6_2,
	lpp_ram_data_out_15_3,
	lpp_ram_data_out_15_0,
	lpp_ram_data_out_15_1,
	lpp_ram_data_out_15_2,
	lpp_ram_data_out_7_3,
	lpp_ram_data_out_7_0,
	lpp_ram_data_out_7_1,
	lpp_ram_data_out_7_2,
	lpp_ram_data_out_9_3,
	lpp_ram_data_out_9_0,
	lpp_ram_data_out_9_1,
	lpp_ram_data_out_9_2,
	lpp_ram_data_out_1_3,
	lpp_ram_data_out_1_0,
	lpp_ram_data_out_1_1,
	lpp_ram_data_out_1_2,
	lpp_ram_data_out_8_3,
	lpp_ram_data_out_8_0,
	lpp_ram_data_out_8_1,
	lpp_ram_data_out_8_2,
	lpp_ram_data_out_0_3,
	lpp_ram_data_out_0_0,
	lpp_ram_data_out_0_1,
	lpp_ram_data_out_0_2,
	global_clock_enable,
	ram_in_reg_2_3,
	ram_in_reg_2_7,
	ram_in_reg_2_1,
	ram_in_reg_2_5,
	ram_in_reg_2_2,
	ram_in_reg_2_0,
	ram_in_reg_2_6,
	ram_in_reg_2_4,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_3_2,
	ram_in_reg_3_0,
	ram_in_reg_3_6,
	ram_in_reg_3_4,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_4_2,
	ram_in_reg_4_0,
	ram_in_reg_4_6,
	ram_in_reg_4_4,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_5_2,
	ram_in_reg_5_0,
	ram_in_reg_5_6,
	ram_in_reg_5_4,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_6_2,
	ram_in_reg_6_0,
	ram_in_reg_6_6,
	ram_in_reg_6_4,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_7_2,
	ram_in_reg_7_0,
	ram_in_reg_7_6,
	ram_in_reg_7_4,
	ram_in_reg_1_3,
	ram_in_reg_1_7,
	ram_in_reg_1_1,
	ram_in_reg_1_5,
	ram_in_reg_1_2,
	ram_in_reg_1_0,
	ram_in_reg_1_6,
	ram_in_reg_1_4,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	ram_in_reg_0_1,
	ram_in_reg_0_5,
	ram_in_reg_0_2,
	ram_in_reg_0_0,
	ram_in_reg_0_6,
	ram_in_reg_0_4,
	clk)/* synthesis synthesis_greybox=1 */;
input 	lpp_ram_data_out_10_3;
input 	lpp_ram_data_out_10_0;
input 	lpp_ram_data_out_10_1;
input 	lpp_ram_data_out_10_2;
input 	tdl_arr_0_4;
input 	tdl_arr_1_4;
input 	lpp_ram_data_out_2_3;
input 	lpp_ram_data_out_2_0;
input 	lpp_ram_data_out_2_1;
input 	lpp_ram_data_out_2_2;
input 	lpp_ram_data_out_11_3;
input 	lpp_ram_data_out_11_0;
input 	lpp_ram_data_out_11_1;
input 	lpp_ram_data_out_11_2;
input 	lpp_ram_data_out_3_3;
input 	lpp_ram_data_out_3_0;
input 	lpp_ram_data_out_3_1;
input 	lpp_ram_data_out_3_2;
input 	lpp_ram_data_out_12_3;
input 	lpp_ram_data_out_12_0;
input 	lpp_ram_data_out_12_1;
input 	lpp_ram_data_out_12_2;
input 	lpp_ram_data_out_4_3;
input 	lpp_ram_data_out_4_0;
input 	lpp_ram_data_out_4_1;
input 	lpp_ram_data_out_4_2;
input 	lpp_ram_data_out_13_3;
input 	lpp_ram_data_out_13_0;
input 	lpp_ram_data_out_13_1;
input 	lpp_ram_data_out_13_2;
input 	lpp_ram_data_out_5_3;
input 	lpp_ram_data_out_5_0;
input 	lpp_ram_data_out_5_1;
input 	lpp_ram_data_out_5_2;
input 	lpp_ram_data_out_14_3;
input 	lpp_ram_data_out_14_0;
input 	lpp_ram_data_out_14_1;
input 	lpp_ram_data_out_14_2;
input 	lpp_ram_data_out_6_3;
input 	lpp_ram_data_out_6_0;
input 	lpp_ram_data_out_6_1;
input 	lpp_ram_data_out_6_2;
input 	lpp_ram_data_out_15_3;
input 	lpp_ram_data_out_15_0;
input 	lpp_ram_data_out_15_1;
input 	lpp_ram_data_out_15_2;
input 	lpp_ram_data_out_7_3;
input 	lpp_ram_data_out_7_0;
input 	lpp_ram_data_out_7_1;
input 	lpp_ram_data_out_7_2;
input 	lpp_ram_data_out_9_3;
input 	lpp_ram_data_out_9_0;
input 	lpp_ram_data_out_9_1;
input 	lpp_ram_data_out_9_2;
input 	lpp_ram_data_out_1_3;
input 	lpp_ram_data_out_1_0;
input 	lpp_ram_data_out_1_1;
input 	lpp_ram_data_out_1_2;
input 	lpp_ram_data_out_8_3;
input 	lpp_ram_data_out_8_0;
input 	lpp_ram_data_out_8_1;
input 	lpp_ram_data_out_8_2;
input 	lpp_ram_data_out_0_3;
input 	lpp_ram_data_out_0_0;
input 	lpp_ram_data_out_0_1;
input 	lpp_ram_data_out_0_2;
input 	global_clock_enable;
output 	ram_in_reg_2_3;
output 	ram_in_reg_2_7;
output 	ram_in_reg_2_1;
output 	ram_in_reg_2_5;
output 	ram_in_reg_2_2;
output 	ram_in_reg_2_0;
output 	ram_in_reg_2_6;
output 	ram_in_reg_2_4;
output 	ram_in_reg_3_3;
output 	ram_in_reg_3_7;
output 	ram_in_reg_3_1;
output 	ram_in_reg_3_5;
output 	ram_in_reg_3_2;
output 	ram_in_reg_3_0;
output 	ram_in_reg_3_6;
output 	ram_in_reg_3_4;
output 	ram_in_reg_4_3;
output 	ram_in_reg_4_7;
output 	ram_in_reg_4_1;
output 	ram_in_reg_4_5;
output 	ram_in_reg_4_2;
output 	ram_in_reg_4_0;
output 	ram_in_reg_4_6;
output 	ram_in_reg_4_4;
output 	ram_in_reg_5_3;
output 	ram_in_reg_5_7;
output 	ram_in_reg_5_1;
output 	ram_in_reg_5_5;
output 	ram_in_reg_5_2;
output 	ram_in_reg_5_0;
output 	ram_in_reg_5_6;
output 	ram_in_reg_5_4;
output 	ram_in_reg_6_3;
output 	ram_in_reg_6_7;
output 	ram_in_reg_6_1;
output 	ram_in_reg_6_5;
output 	ram_in_reg_6_2;
output 	ram_in_reg_6_0;
output 	ram_in_reg_6_6;
output 	ram_in_reg_6_4;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_7;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_5;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_0;
output 	ram_in_reg_7_6;
output 	ram_in_reg_7_4;
output 	ram_in_reg_1_3;
output 	ram_in_reg_1_7;
output 	ram_in_reg_1_1;
output 	ram_in_reg_1_5;
output 	ram_in_reg_1_2;
output 	ram_in_reg_1_0;
output 	ram_in_reg_1_6;
output 	ram_in_reg_1_4;
output 	ram_in_reg_0_3;
output 	ram_in_reg_0_7;
output 	ram_in_reg_0_1;
output 	ram_in_reg_0_5;
output 	ram_in_reg_0_2;
output 	ram_in_reg_0_0;
output 	ram_in_reg_0_6;
output 	ram_in_reg_0_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux5~0_combout ;
wire \Mux45~0_combout ;
wire \Mux5~1_combout ;
wire \Mux45~1_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \Mux4~0_combout ;
wire \Mux44~0_combout ;
wire \Mux4~1_combout ;
wire \Mux44~1_combout ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \Mux3~0_combout ;
wire \Mux43~0_combout ;
wire \Mux3~1_combout ;
wire \Mux43~1_combout ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \Mux2~0_combout ;
wire \Mux42~0_combout ;
wire \Mux2~1_combout ;
wire \Mux42~1_combout ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \Mux1~0_combout ;
wire \Mux41~0_combout ;
wire \Mux1~1_combout ;
wire \Mux41~1_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux0~0_combout ;
wire \Mux40~0_combout ;
wire \Mux0~1_combout ;
wire \Mux40~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux6~0_combout ;
wire \Mux46~0_combout ;
wire \Mux6~1_combout ;
wire \Mux46~1_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \Mux7~0_combout ;
wire \Mux47~0_combout ;
wire \Mux7~1_combout ;
wire \Mux47~1_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux47~2_combout ;
wire \Mux47~3_combout ;


dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\Mux45~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\Mux45~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\Mux5~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux5~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\Mux45~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\Mux45~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\Mux44~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\Mux44~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\Mux4~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux4~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\Mux44~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\Mux44~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\Mux43~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\Mux43~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\Mux3~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux3~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\Mux43~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\Mux43~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\Mux42~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\Mux42~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\Mux2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\Mux2~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\Mux42~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\Mux42~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\Mux41~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\Mux41~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\Mux1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\Mux41~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\Mux41~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\Mux40~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\Mux40~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\Mux0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\Mux0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\Mux40~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\Mux40~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\Mux46~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\Mux46~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux6~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\Mux46~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\Mux46~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\Mux47~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\Mux47~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\Mux7~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux7~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\Mux47~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\Mux47~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!lpp_ram_data_out_10_3),
	.datab(!lpp_ram_data_out_10_0),
	.datac(!lpp_ram_data_out_10_1),
	.datad(!lpp_ram_data_out_10_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux5~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~0 (
	.dataa(!lpp_ram_data_out_2_3),
	.datab(!lpp_ram_data_out_2_0),
	.datac(!lpp_ram_data_out_2_1),
	.datad(!lpp_ram_data_out_2_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~0 .extended_lut = "off";
defparam \Mux45~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~1 (
	.dataa(!lpp_ram_data_out_10_1),
	.datab(!lpp_ram_data_out_10_2),
	.datac(!lpp_ram_data_out_10_3),
	.datad(!lpp_ram_data_out_10_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~1 .extended_lut = "off";
defparam \Mux5~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux5~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~1 (
	.dataa(!lpp_ram_data_out_2_1),
	.datab(!lpp_ram_data_out_2_2),
	.datac(!lpp_ram_data_out_2_3),
	.datad(!lpp_ram_data_out_2_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~1 .extended_lut = "off";
defparam \Mux45~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~2 (
	.dataa(!lpp_ram_data_out_10_2),
	.datab(!lpp_ram_data_out_10_3),
	.datac(!lpp_ram_data_out_10_0),
	.datad(!lpp_ram_data_out_10_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~2 .extended_lut = "off";
defparam \Mux5~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux5~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~3 (
	.dataa(!lpp_ram_data_out_10_0),
	.datab(!lpp_ram_data_out_10_1),
	.datac(!lpp_ram_data_out_10_2),
	.datad(!lpp_ram_data_out_10_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~3 .extended_lut = "off";
defparam \Mux5~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux5~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~2 (
	.dataa(!lpp_ram_data_out_2_2),
	.datab(!lpp_ram_data_out_2_3),
	.datac(!lpp_ram_data_out_2_0),
	.datad(!lpp_ram_data_out_2_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~2 .extended_lut = "off";
defparam \Mux45~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~3 (
	.dataa(!lpp_ram_data_out_2_0),
	.datab(!lpp_ram_data_out_2_1),
	.datac(!lpp_ram_data_out_2_2),
	.datad(!lpp_ram_data_out_2_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~3 .extended_lut = "off";
defparam \Mux45~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!lpp_ram_data_out_11_3),
	.datab(!lpp_ram_data_out_11_0),
	.datac(!lpp_ram_data_out_11_1),
	.datad(!lpp_ram_data_out_11_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~0 (
	.dataa(!lpp_ram_data_out_3_3),
	.datab(!lpp_ram_data_out_3_0),
	.datac(!lpp_ram_data_out_3_1),
	.datad(!lpp_ram_data_out_3_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~0 .extended_lut = "off";
defparam \Mux44~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~1 (
	.dataa(!lpp_ram_data_out_11_1),
	.datab(!lpp_ram_data_out_11_2),
	.datac(!lpp_ram_data_out_11_3),
	.datad(!lpp_ram_data_out_11_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~1 .extended_lut = "off";
defparam \Mux4~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux4~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~1 (
	.dataa(!lpp_ram_data_out_3_1),
	.datab(!lpp_ram_data_out_3_2),
	.datac(!lpp_ram_data_out_3_3),
	.datad(!lpp_ram_data_out_3_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~1 .extended_lut = "off";
defparam \Mux44~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~2 (
	.dataa(!lpp_ram_data_out_11_2),
	.datab(!lpp_ram_data_out_11_3),
	.datac(!lpp_ram_data_out_11_0),
	.datad(!lpp_ram_data_out_11_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~2 .extended_lut = "off";
defparam \Mux4~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux4~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~3 (
	.dataa(!lpp_ram_data_out_11_0),
	.datab(!lpp_ram_data_out_11_1),
	.datac(!lpp_ram_data_out_11_2),
	.datad(!lpp_ram_data_out_11_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~3 .extended_lut = "off";
defparam \Mux4~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux4~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~2 (
	.dataa(!lpp_ram_data_out_3_2),
	.datab(!lpp_ram_data_out_3_3),
	.datac(!lpp_ram_data_out_3_0),
	.datad(!lpp_ram_data_out_3_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~2 .extended_lut = "off";
defparam \Mux44~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~3 (
	.dataa(!lpp_ram_data_out_3_0),
	.datab(!lpp_ram_data_out_3_1),
	.datac(!lpp_ram_data_out_3_2),
	.datad(!lpp_ram_data_out_3_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~3 .extended_lut = "off";
defparam \Mux44~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!lpp_ram_data_out_12_3),
	.datab(!lpp_ram_data_out_12_0),
	.datac(!lpp_ram_data_out_12_1),
	.datad(!lpp_ram_data_out_12_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~0 (
	.dataa(!lpp_ram_data_out_4_3),
	.datab(!lpp_ram_data_out_4_0),
	.datac(!lpp_ram_data_out_4_1),
	.datad(!lpp_ram_data_out_4_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~0 .extended_lut = "off";
defparam \Mux43~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~1 (
	.dataa(!lpp_ram_data_out_12_1),
	.datab(!lpp_ram_data_out_12_2),
	.datac(!lpp_ram_data_out_12_3),
	.datad(!lpp_ram_data_out_12_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~1 .extended_lut = "off";
defparam \Mux3~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux3~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~1 (
	.dataa(!lpp_ram_data_out_4_1),
	.datab(!lpp_ram_data_out_4_2),
	.datac(!lpp_ram_data_out_4_3),
	.datad(!lpp_ram_data_out_4_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~1 .extended_lut = "off";
defparam \Mux43~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~2 (
	.dataa(!lpp_ram_data_out_12_2),
	.datab(!lpp_ram_data_out_12_3),
	.datac(!lpp_ram_data_out_12_0),
	.datad(!lpp_ram_data_out_12_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~2 .extended_lut = "off";
defparam \Mux3~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux3~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~3 (
	.dataa(!lpp_ram_data_out_12_0),
	.datab(!lpp_ram_data_out_12_1),
	.datac(!lpp_ram_data_out_12_2),
	.datad(!lpp_ram_data_out_12_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~3 .extended_lut = "off";
defparam \Mux3~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux3~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~2 (
	.dataa(!lpp_ram_data_out_4_2),
	.datab(!lpp_ram_data_out_4_3),
	.datac(!lpp_ram_data_out_4_0),
	.datad(!lpp_ram_data_out_4_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~2 .extended_lut = "off";
defparam \Mux43~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~3 (
	.dataa(!lpp_ram_data_out_4_0),
	.datab(!lpp_ram_data_out_4_1),
	.datac(!lpp_ram_data_out_4_2),
	.datad(!lpp_ram_data_out_4_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~3 .extended_lut = "off";
defparam \Mux43~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!lpp_ram_data_out_13_3),
	.datab(!lpp_ram_data_out_13_0),
	.datac(!lpp_ram_data_out_13_1),
	.datad(!lpp_ram_data_out_13_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~0 (
	.dataa(!lpp_ram_data_out_5_3),
	.datab(!lpp_ram_data_out_5_0),
	.datac(!lpp_ram_data_out_5_1),
	.datad(!lpp_ram_data_out_5_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~0 .extended_lut = "off";
defparam \Mux42~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~1 (
	.dataa(!lpp_ram_data_out_13_1),
	.datab(!lpp_ram_data_out_13_2),
	.datac(!lpp_ram_data_out_13_3),
	.datad(!lpp_ram_data_out_13_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~1 .extended_lut = "off";
defparam \Mux2~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~1 (
	.dataa(!lpp_ram_data_out_5_1),
	.datab(!lpp_ram_data_out_5_2),
	.datac(!lpp_ram_data_out_5_3),
	.datad(!lpp_ram_data_out_5_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~1 .extended_lut = "off";
defparam \Mux42~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~2 (
	.dataa(!lpp_ram_data_out_13_2),
	.datab(!lpp_ram_data_out_13_3),
	.datac(!lpp_ram_data_out_13_0),
	.datad(!lpp_ram_data_out_13_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~2 .extended_lut = "off";
defparam \Mux2~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~3 (
	.dataa(!lpp_ram_data_out_13_0),
	.datab(!lpp_ram_data_out_13_1),
	.datac(!lpp_ram_data_out_13_2),
	.datad(!lpp_ram_data_out_13_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~3 .extended_lut = "off";
defparam \Mux2~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~2 (
	.dataa(!lpp_ram_data_out_5_2),
	.datab(!lpp_ram_data_out_5_3),
	.datac(!lpp_ram_data_out_5_0),
	.datad(!lpp_ram_data_out_5_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~2 .extended_lut = "off";
defparam \Mux42~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~3 (
	.dataa(!lpp_ram_data_out_5_0),
	.datab(!lpp_ram_data_out_5_1),
	.datac(!lpp_ram_data_out_5_2),
	.datad(!lpp_ram_data_out_5_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~3 .extended_lut = "off";
defparam \Mux42~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!lpp_ram_data_out_14_3),
	.datab(!lpp_ram_data_out_14_0),
	.datac(!lpp_ram_data_out_14_1),
	.datad(!lpp_ram_data_out_14_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~0 (
	.dataa(!lpp_ram_data_out_6_3),
	.datab(!lpp_ram_data_out_6_0),
	.datac(!lpp_ram_data_out_6_1),
	.datad(!lpp_ram_data_out_6_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~0 .extended_lut = "off";
defparam \Mux41~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~1 (
	.dataa(!lpp_ram_data_out_14_1),
	.datab(!lpp_ram_data_out_14_2),
	.datac(!lpp_ram_data_out_14_3),
	.datad(!lpp_ram_data_out_14_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~1 .extended_lut = "off";
defparam \Mux1~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~1 (
	.dataa(!lpp_ram_data_out_6_1),
	.datab(!lpp_ram_data_out_6_2),
	.datac(!lpp_ram_data_out_6_3),
	.datad(!lpp_ram_data_out_6_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~1 .extended_lut = "off";
defparam \Mux41~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~2 (
	.dataa(!lpp_ram_data_out_14_2),
	.datab(!lpp_ram_data_out_14_3),
	.datac(!lpp_ram_data_out_14_0),
	.datad(!lpp_ram_data_out_14_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~2 .extended_lut = "off";
defparam \Mux1~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~3 (
	.dataa(!lpp_ram_data_out_14_0),
	.datab(!lpp_ram_data_out_14_1),
	.datac(!lpp_ram_data_out_14_2),
	.datad(!lpp_ram_data_out_14_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~3 .extended_lut = "off";
defparam \Mux1~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~2 (
	.dataa(!lpp_ram_data_out_6_2),
	.datab(!lpp_ram_data_out_6_3),
	.datac(!lpp_ram_data_out_6_0),
	.datad(!lpp_ram_data_out_6_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~2 .extended_lut = "off";
defparam \Mux41~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~3 (
	.dataa(!lpp_ram_data_out_6_0),
	.datab(!lpp_ram_data_out_6_1),
	.datac(!lpp_ram_data_out_6_2),
	.datad(!lpp_ram_data_out_6_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~3 .extended_lut = "off";
defparam \Mux41~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!lpp_ram_data_out_15_3),
	.datab(!lpp_ram_data_out_15_0),
	.datac(!lpp_ram_data_out_15_1),
	.datad(!lpp_ram_data_out_15_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~0 (
	.dataa(!lpp_ram_data_out_7_3),
	.datab(!lpp_ram_data_out_7_0),
	.datac(!lpp_ram_data_out_7_1),
	.datad(!lpp_ram_data_out_7_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~0 .extended_lut = "off";
defparam \Mux40~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!lpp_ram_data_out_15_1),
	.datab(!lpp_ram_data_out_15_2),
	.datac(!lpp_ram_data_out_15_3),
	.datad(!lpp_ram_data_out_15_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~1 (
	.dataa(!lpp_ram_data_out_7_1),
	.datab(!lpp_ram_data_out_7_2),
	.datac(!lpp_ram_data_out_7_3),
	.datad(!lpp_ram_data_out_7_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~1 .extended_lut = "off";
defparam \Mux40~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~2 (
	.dataa(!lpp_ram_data_out_15_2),
	.datab(!lpp_ram_data_out_15_3),
	.datac(!lpp_ram_data_out_15_0),
	.datad(!lpp_ram_data_out_15_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~2 .extended_lut = "off";
defparam \Mux0~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~3 (
	.dataa(!lpp_ram_data_out_15_0),
	.datab(!lpp_ram_data_out_15_1),
	.datac(!lpp_ram_data_out_15_2),
	.datad(!lpp_ram_data_out_15_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~3 .extended_lut = "off";
defparam \Mux0~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~2 (
	.dataa(!lpp_ram_data_out_7_2),
	.datab(!lpp_ram_data_out_7_3),
	.datac(!lpp_ram_data_out_7_0),
	.datad(!lpp_ram_data_out_7_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~2 .extended_lut = "off";
defparam \Mux40~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~3 (
	.dataa(!lpp_ram_data_out_7_0),
	.datab(!lpp_ram_data_out_7_1),
	.datac(!lpp_ram_data_out_7_2),
	.datad(!lpp_ram_data_out_7_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~3 .extended_lut = "off";
defparam \Mux40~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!lpp_ram_data_out_9_3),
	.datab(!lpp_ram_data_out_9_0),
	.datac(!lpp_ram_data_out_9_1),
	.datad(!lpp_ram_data_out_9_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~0 (
	.dataa(!lpp_ram_data_out_1_3),
	.datab(!lpp_ram_data_out_1_0),
	.datac(!lpp_ram_data_out_1_1),
	.datad(!lpp_ram_data_out_1_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~0 .extended_lut = "off";
defparam \Mux46~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~1 (
	.dataa(!lpp_ram_data_out_9_1),
	.datab(!lpp_ram_data_out_9_2),
	.datac(!lpp_ram_data_out_9_3),
	.datad(!lpp_ram_data_out_9_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~1 .extended_lut = "off";
defparam \Mux6~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~1 (
	.dataa(!lpp_ram_data_out_1_1),
	.datab(!lpp_ram_data_out_1_2),
	.datac(!lpp_ram_data_out_1_3),
	.datad(!lpp_ram_data_out_1_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~1 .extended_lut = "off";
defparam \Mux46~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~2 (
	.dataa(!lpp_ram_data_out_9_2),
	.datab(!lpp_ram_data_out_9_3),
	.datac(!lpp_ram_data_out_9_0),
	.datad(!lpp_ram_data_out_9_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~2 .extended_lut = "off";
defparam \Mux6~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~3 (
	.dataa(!lpp_ram_data_out_9_0),
	.datab(!lpp_ram_data_out_9_1),
	.datac(!lpp_ram_data_out_9_2),
	.datad(!lpp_ram_data_out_9_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~3 .extended_lut = "off";
defparam \Mux6~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~2 (
	.dataa(!lpp_ram_data_out_1_2),
	.datab(!lpp_ram_data_out_1_3),
	.datac(!lpp_ram_data_out_1_0),
	.datad(!lpp_ram_data_out_1_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~2 .extended_lut = "off";
defparam \Mux46~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~3 (
	.dataa(!lpp_ram_data_out_1_0),
	.datab(!lpp_ram_data_out_1_1),
	.datac(!lpp_ram_data_out_1_2),
	.datad(!lpp_ram_data_out_1_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~3 .extended_lut = "off";
defparam \Mux46~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!lpp_ram_data_out_8_3),
	.datab(!lpp_ram_data_out_8_0),
	.datac(!lpp_ram_data_out_8_1),
	.datad(!lpp_ram_data_out_8_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~0 (
	.dataa(!lpp_ram_data_out_0_3),
	.datab(!lpp_ram_data_out_0_0),
	.datac(!lpp_ram_data_out_0_1),
	.datad(!lpp_ram_data_out_0_2),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~0 .extended_lut = "off";
defparam \Mux47~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~1 (
	.dataa(!lpp_ram_data_out_8_1),
	.datab(!lpp_ram_data_out_8_2),
	.datac(!lpp_ram_data_out_8_3),
	.datad(!lpp_ram_data_out_8_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~1 .extended_lut = "off";
defparam \Mux7~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux7~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~1 (
	.dataa(!lpp_ram_data_out_0_1),
	.datab(!lpp_ram_data_out_0_2),
	.datac(!lpp_ram_data_out_0_3),
	.datad(!lpp_ram_data_out_0_0),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~1 .extended_lut = "off";
defparam \Mux47~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~2 (
	.dataa(!lpp_ram_data_out_8_2),
	.datab(!lpp_ram_data_out_8_3),
	.datac(!lpp_ram_data_out_8_0),
	.datad(!lpp_ram_data_out_8_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~2 .extended_lut = "off";
defparam \Mux7~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux7~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~3 (
	.dataa(!lpp_ram_data_out_8_0),
	.datab(!lpp_ram_data_out_8_1),
	.datac(!lpp_ram_data_out_8_2),
	.datad(!lpp_ram_data_out_8_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~3 .extended_lut = "off";
defparam \Mux7~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux7~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~2 (
	.dataa(!lpp_ram_data_out_0_2),
	.datab(!lpp_ram_data_out_0_3),
	.datac(!lpp_ram_data_out_0_0),
	.datad(!lpp_ram_data_out_0_1),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~2 .extended_lut = "off";
defparam \Mux47~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~3 (
	.dataa(!lpp_ram_data_out_0_0),
	.datab(!lpp_ram_data_out_0_1),
	.datac(!lpp_ram_data_out_0_2),
	.datad(!lpp_ram_data_out_0_3),
	.datae(!tdl_arr_0_4),
	.dataf(!tdl_arr_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~3 .extended_lut = "off";
defparam \Mux47~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~3 .shared_arith = "off";

endmodule

module IFFT_asj_fft_cxb_data_r_1 (
	global_clock_enable,
	ram_in_reg_6_1,
	ram_in_reg_5_1,
	ram_in_reg_2_1,
	ram_in_reg_3_1,
	ram_in_reg_4_1,
	ram_in_reg_6_3,
	ram_in_reg_5_3,
	ram_in_reg_2_3,
	ram_in_reg_3_3,
	ram_in_reg_4_3,
	ram_in_reg_6_0,
	ram_in_reg_5_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_6_2,
	ram_in_reg_5_2,
	ram_in_reg_2_2,
	ram_in_reg_3_2,
	ram_in_reg_4_2,
	ram_in_reg_7_1,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_2,
	ram_in_reg_7_5,
	ram_in_reg_6_5,
	ram_in_reg_3_5,
	ram_in_reg_4_5,
	ram_in_reg_5_5,
	ram_in_reg_7_7,
	ram_in_reg_6_7,
	ram_in_reg_3_7,
	ram_in_reg_4_7,
	ram_in_reg_5_7,
	ram_in_reg_7_4,
	ram_in_reg_6_4,
	ram_in_reg_3_4,
	ram_in_reg_4_4,
	ram_in_reg_5_4,
	ram_in_reg_7_6,
	ram_in_reg_6_6,
	ram_in_reg_3_6,
	ram_in_reg_4_6,
	ram_in_reg_5_6,
	ram_in_reg_2_5,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_6,
	ram_in_reg_0_2,
	ram_in_reg_1_2,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_0_7,
	ram_in_reg_1_7,
	ram_in_reg_0_5,
	ram_in_reg_1_5,
	ram_in_reg_0_3,
	ram_in_reg_1_3,
	ram_in_reg_0_1,
	ram_in_reg_1_1,
	ram_in_reg_0_6,
	ram_in_reg_1_6,
	ram_in_reg_0_4,
	ram_in_reg_1_4,
	ram_data_out1_14,
	ram_data_out2_14,
	ram_data_out3_14,
	ram_data_out0_14,
	sw_r_tdl_0_4,
	sw_r_tdl_1_4,
	ram_data_out1_13,
	ram_data_out2_13,
	ram_data_out3_13,
	ram_data_out0_13,
	ram_data_out1_10,
	ram_data_out2_10,
	ram_data_out3_10,
	ram_data_out0_10,
	ram_data_out1_11,
	ram_data_out2_11,
	ram_data_out3_11,
	ram_data_out0_11,
	ram_data_out1_12,
	ram_data_out2_12,
	ram_data_out3_12,
	ram_data_out0_12,
	ram_data_out1_15,
	ram_data_out2_15,
	ram_data_out3_15,
	ram_data_out0_15,
	ram_data_out1_7,
	ram_data_out2_7,
	ram_data_out3_7,
	ram_data_out0_7,
	ram_data_out1_6,
	ram_data_out2_6,
	ram_data_out3_6,
	ram_data_out0_6,
	ram_data_out1_3,
	ram_data_out2_3,
	ram_data_out3_3,
	ram_data_out0_3,
	ram_data_out1_4,
	ram_data_out2_4,
	ram_data_out3_4,
	ram_data_out0_4,
	ram_data_out1_5,
	ram_data_out2_5,
	ram_data_out3_5,
	ram_data_out0_5,
	ram_data_out1_2,
	ram_data_out2_2,
	ram_data_out3_2,
	ram_data_out0_2,
	ram_data_out2_8,
	ram_data_out3_8,
	ram_data_out0_8,
	ram_data_out1_8,
	ram_data_out2_9,
	ram_data_out3_9,
	ram_data_out0_9,
	ram_data_out1_9,
	ram_data_out3_0,
	ram_data_out0_0,
	ram_data_out1_0,
	ram_data_out2_0,
	ram_data_out3_1,
	ram_data_out0_1,
	ram_data_out1_1,
	ram_data_out2_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	ram_in_reg_6_1;
output 	ram_in_reg_5_1;
output 	ram_in_reg_2_1;
output 	ram_in_reg_3_1;
output 	ram_in_reg_4_1;
output 	ram_in_reg_6_3;
output 	ram_in_reg_5_3;
output 	ram_in_reg_2_3;
output 	ram_in_reg_3_3;
output 	ram_in_reg_4_3;
output 	ram_in_reg_6_0;
output 	ram_in_reg_5_0;
output 	ram_in_reg_2_0;
output 	ram_in_reg_3_0;
output 	ram_in_reg_4_0;
output 	ram_in_reg_6_2;
output 	ram_in_reg_5_2;
output 	ram_in_reg_2_2;
output 	ram_in_reg_3_2;
output 	ram_in_reg_4_2;
output 	ram_in_reg_7_1;
output 	ram_in_reg_7_3;
output 	ram_in_reg_7_0;
output 	ram_in_reg_7_2;
output 	ram_in_reg_7_5;
output 	ram_in_reg_6_5;
output 	ram_in_reg_3_5;
output 	ram_in_reg_4_5;
output 	ram_in_reg_5_5;
output 	ram_in_reg_7_7;
output 	ram_in_reg_6_7;
output 	ram_in_reg_3_7;
output 	ram_in_reg_4_7;
output 	ram_in_reg_5_7;
output 	ram_in_reg_7_4;
output 	ram_in_reg_6_4;
output 	ram_in_reg_3_4;
output 	ram_in_reg_4_4;
output 	ram_in_reg_5_4;
output 	ram_in_reg_7_6;
output 	ram_in_reg_6_6;
output 	ram_in_reg_3_6;
output 	ram_in_reg_4_6;
output 	ram_in_reg_5_6;
output 	ram_in_reg_2_5;
output 	ram_in_reg_2_7;
output 	ram_in_reg_2_4;
output 	ram_in_reg_2_6;
output 	ram_in_reg_0_2;
output 	ram_in_reg_1_2;
output 	ram_in_reg_0_0;
output 	ram_in_reg_1_0;
output 	ram_in_reg_0_7;
output 	ram_in_reg_1_7;
output 	ram_in_reg_0_5;
output 	ram_in_reg_1_5;
output 	ram_in_reg_0_3;
output 	ram_in_reg_1_3;
output 	ram_in_reg_0_1;
output 	ram_in_reg_1_1;
output 	ram_in_reg_0_6;
output 	ram_in_reg_1_6;
output 	ram_in_reg_0_4;
output 	ram_in_reg_1_4;
input 	ram_data_out1_14;
input 	ram_data_out2_14;
input 	ram_data_out3_14;
input 	ram_data_out0_14;
input 	sw_r_tdl_0_4;
input 	sw_r_tdl_1_4;
input 	ram_data_out1_13;
input 	ram_data_out2_13;
input 	ram_data_out3_13;
input 	ram_data_out0_13;
input 	ram_data_out1_10;
input 	ram_data_out2_10;
input 	ram_data_out3_10;
input 	ram_data_out0_10;
input 	ram_data_out1_11;
input 	ram_data_out2_11;
input 	ram_data_out3_11;
input 	ram_data_out0_11;
input 	ram_data_out1_12;
input 	ram_data_out2_12;
input 	ram_data_out3_12;
input 	ram_data_out0_12;
input 	ram_data_out1_15;
input 	ram_data_out2_15;
input 	ram_data_out3_15;
input 	ram_data_out0_15;
input 	ram_data_out1_7;
input 	ram_data_out2_7;
input 	ram_data_out3_7;
input 	ram_data_out0_7;
input 	ram_data_out1_6;
input 	ram_data_out2_6;
input 	ram_data_out3_6;
input 	ram_data_out0_6;
input 	ram_data_out1_3;
input 	ram_data_out2_3;
input 	ram_data_out3_3;
input 	ram_data_out0_3;
input 	ram_data_out1_4;
input 	ram_data_out2_4;
input 	ram_data_out3_4;
input 	ram_data_out0_4;
input 	ram_data_out1_5;
input 	ram_data_out2_5;
input 	ram_data_out3_5;
input 	ram_data_out0_5;
input 	ram_data_out1_2;
input 	ram_data_out2_2;
input 	ram_data_out3_2;
input 	ram_data_out0_2;
input 	ram_data_out2_8;
input 	ram_data_out3_8;
input 	ram_data_out0_8;
input 	ram_data_out1_8;
input 	ram_data_out2_9;
input 	ram_data_out3_9;
input 	ram_data_out0_9;
input 	ram_data_out1_9;
input 	ram_data_out3_0;
input 	ram_data_out0_0;
input 	ram_data_out1_0;
input 	ram_data_out2_0;
input 	ram_data_out3_1;
input 	ram_data_out0_1;
input 	ram_data_out1_1;
input 	ram_data_out2_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux9~0_combout ;
wire \Mux10~0_combout ;
wire \Mux13~0_combout ;
wire \Mux12~0_combout ;
wire \Mux11~0_combout ;
wire \Mux9~1_combout ;
wire \Mux10~1_combout ;
wire \Mux13~1_combout ;
wire \Mux12~1_combout ;
wire \Mux11~1_combout ;
wire \Mux9~2_combout ;
wire \Mux10~2_combout ;
wire \Mux13~2_combout ;
wire \Mux12~2_combout ;
wire \Mux11~2_combout ;
wire \Mux9~3_combout ;
wire \Mux10~3_combout ;
wire \Mux13~3_combout ;
wire \Mux12~3_combout ;
wire \Mux11~3_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux40~0_combout ;
wire \Mux41~0_combout ;
wire \Mux44~0_combout ;
wire \Mux43~0_combout ;
wire \Mux42~0_combout ;
wire \Mux40~1_combout ;
wire \Mux41~1_combout ;
wire \Mux44~1_combout ;
wire \Mux43~1_combout ;
wire \Mux42~1_combout ;
wire \Mux40~2_combout ;
wire \Mux41~2_combout ;
wire \Mux44~2_combout ;
wire \Mux43~2_combout ;
wire \Mux42~2_combout ;
wire \Mux40~3_combout ;
wire \Mux41~3_combout ;
wire \Mux44~3_combout ;
wire \Mux43~3_combout ;
wire \Mux42~3_combout ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \Mux15~0_combout ;
wire \Mux14~0_combout ;
wire \Mux15~1_combout ;
wire \Mux14~1_combout ;
wire \Mux47~0_combout ;
wire \Mux46~0_combout ;
wire \Mux47~1_combout ;
wire \Mux46~1_combout ;
wire \Mux15~2_combout ;
wire \Mux14~2_combout ;
wire \Mux15~3_combout ;
wire \Mux14~3_combout ;
wire \Mux47~2_combout ;
wire \Mux46~2_combout ;
wire \Mux47~3_combout ;
wire \Mux46~3_combout ;


dffeas \ram_in_reg[1][6] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_1),
	.prn(vcc));
defparam \ram_in_reg[1][6] .is_wysiwyg = "true";
defparam \ram_in_reg[1][6] .power_up = "low";

dffeas \ram_in_reg[1][5] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_1),
	.prn(vcc));
defparam \ram_in_reg[1][5] .is_wysiwyg = "true";
defparam \ram_in_reg[1][5] .power_up = "low";

dffeas \ram_in_reg[1][2] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_1),
	.prn(vcc));
defparam \ram_in_reg[1][2] .is_wysiwyg = "true";
defparam \ram_in_reg[1][2] .power_up = "low";

dffeas \ram_in_reg[1][3] (
	.clk(clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_1),
	.prn(vcc));
defparam \ram_in_reg[1][3] .is_wysiwyg = "true";
defparam \ram_in_reg[1][3] .power_up = "low";

dffeas \ram_in_reg[1][4] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_1),
	.prn(vcc));
defparam \ram_in_reg[1][4] .is_wysiwyg = "true";
defparam \ram_in_reg[1][4] .power_up = "low";

dffeas \ram_in_reg[3][6] (
	.clk(clk),
	.d(\Mux9~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_3),
	.prn(vcc));
defparam \ram_in_reg[3][6] .is_wysiwyg = "true";
defparam \ram_in_reg[3][6] .power_up = "low";

dffeas \ram_in_reg[3][5] (
	.clk(clk),
	.d(\Mux10~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_3),
	.prn(vcc));
defparam \ram_in_reg[3][5] .is_wysiwyg = "true";
defparam \ram_in_reg[3][5] .power_up = "low";

dffeas \ram_in_reg[3][2] (
	.clk(clk),
	.d(\Mux13~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_3),
	.prn(vcc));
defparam \ram_in_reg[3][2] .is_wysiwyg = "true";
defparam \ram_in_reg[3][2] .power_up = "low";

dffeas \ram_in_reg[3][3] (
	.clk(clk),
	.d(\Mux12~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_3),
	.prn(vcc));
defparam \ram_in_reg[3][3] .is_wysiwyg = "true";
defparam \ram_in_reg[3][3] .power_up = "low";

dffeas \ram_in_reg[3][4] (
	.clk(clk),
	.d(\Mux11~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_3),
	.prn(vcc));
defparam \ram_in_reg[3][4] .is_wysiwyg = "true";
defparam \ram_in_reg[3][4] .power_up = "low";

dffeas \ram_in_reg[0][6] (
	.clk(clk),
	.d(\Mux9~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_0),
	.prn(vcc));
defparam \ram_in_reg[0][6] .is_wysiwyg = "true";
defparam \ram_in_reg[0][6] .power_up = "low";

dffeas \ram_in_reg[0][5] (
	.clk(clk),
	.d(\Mux10~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_0),
	.prn(vcc));
defparam \ram_in_reg[0][5] .is_wysiwyg = "true";
defparam \ram_in_reg[0][5] .power_up = "low";

dffeas \ram_in_reg[0][2] (
	.clk(clk),
	.d(\Mux13~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_0),
	.prn(vcc));
defparam \ram_in_reg[0][2] .is_wysiwyg = "true";
defparam \ram_in_reg[0][2] .power_up = "low";

dffeas \ram_in_reg[0][3] (
	.clk(clk),
	.d(\Mux12~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_0),
	.prn(vcc));
defparam \ram_in_reg[0][3] .is_wysiwyg = "true";
defparam \ram_in_reg[0][3] .power_up = "low";

dffeas \ram_in_reg[0][4] (
	.clk(clk),
	.d(\Mux11~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_0),
	.prn(vcc));
defparam \ram_in_reg[0][4] .is_wysiwyg = "true";
defparam \ram_in_reg[0][4] .power_up = "low";

dffeas \ram_in_reg[2][6] (
	.clk(clk),
	.d(\Mux9~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_2),
	.prn(vcc));
defparam \ram_in_reg[2][6] .is_wysiwyg = "true";
defparam \ram_in_reg[2][6] .power_up = "low";

dffeas \ram_in_reg[2][5] (
	.clk(clk),
	.d(\Mux10~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_2),
	.prn(vcc));
defparam \ram_in_reg[2][5] .is_wysiwyg = "true";
defparam \ram_in_reg[2][5] .power_up = "low";

dffeas \ram_in_reg[2][2] (
	.clk(clk),
	.d(\Mux13~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_2),
	.prn(vcc));
defparam \ram_in_reg[2][2] .is_wysiwyg = "true";
defparam \ram_in_reg[2][2] .power_up = "low";

dffeas \ram_in_reg[2][3] (
	.clk(clk),
	.d(\Mux12~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_2),
	.prn(vcc));
defparam \ram_in_reg[2][3] .is_wysiwyg = "true";
defparam \ram_in_reg[2][3] .power_up = "low";

dffeas \ram_in_reg[2][4] (
	.clk(clk),
	.d(\Mux11~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_2),
	.prn(vcc));
defparam \ram_in_reg[2][4] .is_wysiwyg = "true";
defparam \ram_in_reg[2][4] .power_up = "low";

dffeas \ram_in_reg[1][7] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_1),
	.prn(vcc));
defparam \ram_in_reg[1][7] .is_wysiwyg = "true";
defparam \ram_in_reg[1][7] .power_up = "low";

dffeas \ram_in_reg[3][7] (
	.clk(clk),
	.d(\Mux8~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_3),
	.prn(vcc));
defparam \ram_in_reg[3][7] .is_wysiwyg = "true";
defparam \ram_in_reg[3][7] .power_up = "low";

dffeas \ram_in_reg[0][7] (
	.clk(clk),
	.d(\Mux8~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_0),
	.prn(vcc));
defparam \ram_in_reg[0][7] .is_wysiwyg = "true";
defparam \ram_in_reg[0][7] .power_up = "low";

dffeas \ram_in_reg[2][7] (
	.clk(clk),
	.d(\Mux8~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_2),
	.prn(vcc));
defparam \ram_in_reg[2][7] .is_wysiwyg = "true";
defparam \ram_in_reg[2][7] .power_up = "low";

dffeas \ram_in_reg[5][7] (
	.clk(clk),
	.d(\Mux40~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_5),
	.prn(vcc));
defparam \ram_in_reg[5][7] .is_wysiwyg = "true";
defparam \ram_in_reg[5][7] .power_up = "low";

dffeas \ram_in_reg[5][6] (
	.clk(clk),
	.d(\Mux41~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_5),
	.prn(vcc));
defparam \ram_in_reg[5][6] .is_wysiwyg = "true";
defparam \ram_in_reg[5][6] .power_up = "low";

dffeas \ram_in_reg[5][3] (
	.clk(clk),
	.d(\Mux44~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_5),
	.prn(vcc));
defparam \ram_in_reg[5][3] .is_wysiwyg = "true";
defparam \ram_in_reg[5][3] .power_up = "low";

dffeas \ram_in_reg[5][4] (
	.clk(clk),
	.d(\Mux43~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_5),
	.prn(vcc));
defparam \ram_in_reg[5][4] .is_wysiwyg = "true";
defparam \ram_in_reg[5][4] .power_up = "low";

dffeas \ram_in_reg[5][5] (
	.clk(clk),
	.d(\Mux42~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_5),
	.prn(vcc));
defparam \ram_in_reg[5][5] .is_wysiwyg = "true";
defparam \ram_in_reg[5][5] .power_up = "low";

dffeas \ram_in_reg[7][7] (
	.clk(clk),
	.d(\Mux40~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_7),
	.prn(vcc));
defparam \ram_in_reg[7][7] .is_wysiwyg = "true";
defparam \ram_in_reg[7][7] .power_up = "low";

dffeas \ram_in_reg[7][6] (
	.clk(clk),
	.d(\Mux41~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_7),
	.prn(vcc));
defparam \ram_in_reg[7][6] .is_wysiwyg = "true";
defparam \ram_in_reg[7][6] .power_up = "low";

dffeas \ram_in_reg[7][3] (
	.clk(clk),
	.d(\Mux44~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_7),
	.prn(vcc));
defparam \ram_in_reg[7][3] .is_wysiwyg = "true";
defparam \ram_in_reg[7][3] .power_up = "low";

dffeas \ram_in_reg[7][4] (
	.clk(clk),
	.d(\Mux43~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_7),
	.prn(vcc));
defparam \ram_in_reg[7][4] .is_wysiwyg = "true";
defparam \ram_in_reg[7][4] .power_up = "low";

dffeas \ram_in_reg[7][5] (
	.clk(clk),
	.d(\Mux42~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_7),
	.prn(vcc));
defparam \ram_in_reg[7][5] .is_wysiwyg = "true";
defparam \ram_in_reg[7][5] .power_up = "low";

dffeas \ram_in_reg[4][7] (
	.clk(clk),
	.d(\Mux40~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_4),
	.prn(vcc));
defparam \ram_in_reg[4][7] .is_wysiwyg = "true";
defparam \ram_in_reg[4][7] .power_up = "low";

dffeas \ram_in_reg[4][6] (
	.clk(clk),
	.d(\Mux41~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_4),
	.prn(vcc));
defparam \ram_in_reg[4][6] .is_wysiwyg = "true";
defparam \ram_in_reg[4][6] .power_up = "low";

dffeas \ram_in_reg[4][3] (
	.clk(clk),
	.d(\Mux44~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_4),
	.prn(vcc));
defparam \ram_in_reg[4][3] .is_wysiwyg = "true";
defparam \ram_in_reg[4][3] .power_up = "low";

dffeas \ram_in_reg[4][4] (
	.clk(clk),
	.d(\Mux43~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_4),
	.prn(vcc));
defparam \ram_in_reg[4][4] .is_wysiwyg = "true";
defparam \ram_in_reg[4][4] .power_up = "low";

dffeas \ram_in_reg[4][5] (
	.clk(clk),
	.d(\Mux42~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_4),
	.prn(vcc));
defparam \ram_in_reg[4][5] .is_wysiwyg = "true";
defparam \ram_in_reg[4][5] .power_up = "low";

dffeas \ram_in_reg[6][7] (
	.clk(clk),
	.d(\Mux40~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_7_6),
	.prn(vcc));
defparam \ram_in_reg[6][7] .is_wysiwyg = "true";
defparam \ram_in_reg[6][7] .power_up = "low";

dffeas \ram_in_reg[6][6] (
	.clk(clk),
	.d(\Mux41~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_6_6),
	.prn(vcc));
defparam \ram_in_reg[6][6] .is_wysiwyg = "true";
defparam \ram_in_reg[6][6] .power_up = "low";

dffeas \ram_in_reg[6][3] (
	.clk(clk),
	.d(\Mux44~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_3_6),
	.prn(vcc));
defparam \ram_in_reg[6][3] .is_wysiwyg = "true";
defparam \ram_in_reg[6][3] .power_up = "low";

dffeas \ram_in_reg[6][4] (
	.clk(clk),
	.d(\Mux43~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_4_6),
	.prn(vcc));
defparam \ram_in_reg[6][4] .is_wysiwyg = "true";
defparam \ram_in_reg[6][4] .power_up = "low";

dffeas \ram_in_reg[6][5] (
	.clk(clk),
	.d(\Mux42~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_5_6),
	.prn(vcc));
defparam \ram_in_reg[6][5] .is_wysiwyg = "true";
defparam \ram_in_reg[6][5] .power_up = "low";

dffeas \ram_in_reg[5][2] (
	.clk(clk),
	.d(\Mux45~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_5),
	.prn(vcc));
defparam \ram_in_reg[5][2] .is_wysiwyg = "true";
defparam \ram_in_reg[5][2] .power_up = "low";

dffeas \ram_in_reg[7][2] (
	.clk(clk),
	.d(\Mux45~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_7),
	.prn(vcc));
defparam \ram_in_reg[7][2] .is_wysiwyg = "true";
defparam \ram_in_reg[7][2] .power_up = "low";

dffeas \ram_in_reg[4][2] (
	.clk(clk),
	.d(\Mux45~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_4),
	.prn(vcc));
defparam \ram_in_reg[4][2] .is_wysiwyg = "true";
defparam \ram_in_reg[4][2] .power_up = "low";

dffeas \ram_in_reg[6][2] (
	.clk(clk),
	.d(\Mux45~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_2_6),
	.prn(vcc));
defparam \ram_in_reg[6][2] .is_wysiwyg = "true";
defparam \ram_in_reg[6][2] .power_up = "low";

dffeas \ram_in_reg[2][0] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_2),
	.prn(vcc));
defparam \ram_in_reg[2][0] .is_wysiwyg = "true";
defparam \ram_in_reg[2][0] .power_up = "low";

dffeas \ram_in_reg[2][1] (
	.clk(clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_2),
	.prn(vcc));
defparam \ram_in_reg[2][1] .is_wysiwyg = "true";
defparam \ram_in_reg[2][1] .power_up = "low";

dffeas \ram_in_reg[0][0] (
	.clk(clk),
	.d(\Mux15~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_0),
	.prn(vcc));
defparam \ram_in_reg[0][0] .is_wysiwyg = "true";
defparam \ram_in_reg[0][0] .power_up = "low";

dffeas \ram_in_reg[0][1] (
	.clk(clk),
	.d(\Mux14~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_0),
	.prn(vcc));
defparam \ram_in_reg[0][1] .is_wysiwyg = "true";
defparam \ram_in_reg[0][1] .power_up = "low";

dffeas \ram_in_reg[7][0] (
	.clk(clk),
	.d(\Mux47~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_7),
	.prn(vcc));
defparam \ram_in_reg[7][0] .is_wysiwyg = "true";
defparam \ram_in_reg[7][0] .power_up = "low";

dffeas \ram_in_reg[7][1] (
	.clk(clk),
	.d(\Mux46~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_7),
	.prn(vcc));
defparam \ram_in_reg[7][1] .is_wysiwyg = "true";
defparam \ram_in_reg[7][1] .power_up = "low";

dffeas \ram_in_reg[5][0] (
	.clk(clk),
	.d(\Mux47~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_5),
	.prn(vcc));
defparam \ram_in_reg[5][0] .is_wysiwyg = "true";
defparam \ram_in_reg[5][0] .power_up = "low";

dffeas \ram_in_reg[5][1] (
	.clk(clk),
	.d(\Mux46~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_5),
	.prn(vcc));
defparam \ram_in_reg[5][1] .is_wysiwyg = "true";
defparam \ram_in_reg[5][1] .power_up = "low";

dffeas \ram_in_reg[3][0] (
	.clk(clk),
	.d(\Mux15~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_3),
	.prn(vcc));
defparam \ram_in_reg[3][0] .is_wysiwyg = "true";
defparam \ram_in_reg[3][0] .power_up = "low";

dffeas \ram_in_reg[3][1] (
	.clk(clk),
	.d(\Mux14~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_3),
	.prn(vcc));
defparam \ram_in_reg[3][1] .is_wysiwyg = "true";
defparam \ram_in_reg[3][1] .power_up = "low";

dffeas \ram_in_reg[1][0] (
	.clk(clk),
	.d(\Mux15~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_1),
	.prn(vcc));
defparam \ram_in_reg[1][0] .is_wysiwyg = "true";
defparam \ram_in_reg[1][0] .power_up = "low";

dffeas \ram_in_reg[1][1] (
	.clk(clk),
	.d(\Mux14~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_1),
	.prn(vcc));
defparam \ram_in_reg[1][1] .is_wysiwyg = "true";
defparam \ram_in_reg[1][1] .power_up = "low";

dffeas \ram_in_reg[6][0] (
	.clk(clk),
	.d(\Mux47~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_6),
	.prn(vcc));
defparam \ram_in_reg[6][0] .is_wysiwyg = "true";
defparam \ram_in_reg[6][0] .power_up = "low";

dffeas \ram_in_reg[6][1] (
	.clk(clk),
	.d(\Mux46~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_6),
	.prn(vcc));
defparam \ram_in_reg[6][1] .is_wysiwyg = "true";
defparam \ram_in_reg[6][1] .power_up = "low";

dffeas \ram_in_reg[4][0] (
	.clk(clk),
	.d(\Mux47~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_0_4),
	.prn(vcc));
defparam \ram_in_reg[4][0] .is_wysiwyg = "true";
defparam \ram_in_reg[4][0] .power_up = "low";

dffeas \ram_in_reg[4][1] (
	.clk(clk),
	.d(\Mux46~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(ram_in_reg_1_4),
	.prn(vcc));
defparam \ram_in_reg[4][1] .is_wysiwyg = "true";
defparam \ram_in_reg[4][1] .power_up = "low";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!ram_data_out1_14),
	.datab(!ram_data_out2_14),
	.datac(!ram_data_out3_14),
	.datad(!ram_data_out0_14),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!ram_data_out1_13),
	.datab(!ram_data_out2_13),
	.datac(!ram_data_out3_13),
	.datad(!ram_data_out0_13),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~0 (
	.dataa(!ram_data_out1_10),
	.datab(!ram_data_out2_10),
	.datac(!ram_data_out3_10),
	.datad(!ram_data_out0_10),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "off";
defparam \Mux13~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux13~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~0 (
	.dataa(!ram_data_out1_11),
	.datab(!ram_data_out2_11),
	.datac(!ram_data_out3_11),
	.datad(!ram_data_out0_11),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "off";
defparam \Mux12~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux12~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!ram_data_out1_12),
	.datab(!ram_data_out2_12),
	.datac(!ram_data_out3_12),
	.datad(!ram_data_out0_12),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~1 (
	.dataa(!ram_data_out3_14),
	.datab(!ram_data_out0_14),
	.datac(!ram_data_out1_14),
	.datad(!ram_data_out2_14),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~1 .extended_lut = "off";
defparam \Mux9~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~1 (
	.dataa(!ram_data_out3_13),
	.datab(!ram_data_out0_13),
	.datac(!ram_data_out1_13),
	.datad(!ram_data_out2_13),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~1 .extended_lut = "off";
defparam \Mux10~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~1 (
	.dataa(!ram_data_out3_10),
	.datab(!ram_data_out0_10),
	.datac(!ram_data_out1_10),
	.datad(!ram_data_out2_10),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~1 .extended_lut = "off";
defparam \Mux13~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux13~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~1 (
	.dataa(!ram_data_out3_11),
	.datab(!ram_data_out0_11),
	.datac(!ram_data_out1_11),
	.datad(!ram_data_out2_11),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~1 .extended_lut = "off";
defparam \Mux12~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux12~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~1 (
	.dataa(!ram_data_out3_12),
	.datab(!ram_data_out0_12),
	.datac(!ram_data_out1_12),
	.datad(!ram_data_out2_12),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~1 .extended_lut = "off";
defparam \Mux11~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux11~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~2 (
	.dataa(!ram_data_out0_14),
	.datab(!ram_data_out1_14),
	.datac(!ram_data_out2_14),
	.datad(!ram_data_out3_14),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~2 .extended_lut = "off";
defparam \Mux9~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~2 (
	.dataa(!ram_data_out0_13),
	.datab(!ram_data_out1_13),
	.datac(!ram_data_out2_13),
	.datad(!ram_data_out3_13),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~2 .extended_lut = "off";
defparam \Mux10~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~2 (
	.dataa(!ram_data_out0_10),
	.datab(!ram_data_out1_10),
	.datac(!ram_data_out2_10),
	.datad(!ram_data_out3_10),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~2 .extended_lut = "off";
defparam \Mux13~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux13~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~2 (
	.dataa(!ram_data_out0_11),
	.datab(!ram_data_out1_11),
	.datac(!ram_data_out2_11),
	.datad(!ram_data_out3_11),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~2 .extended_lut = "off";
defparam \Mux12~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux12~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~2 (
	.dataa(!ram_data_out0_12),
	.datab(!ram_data_out1_12),
	.datac(!ram_data_out2_12),
	.datad(!ram_data_out3_12),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~2 .extended_lut = "off";
defparam \Mux11~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux11~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~3 (
	.dataa(!ram_data_out2_14),
	.datab(!ram_data_out3_14),
	.datac(!ram_data_out0_14),
	.datad(!ram_data_out1_14),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~3 .extended_lut = "off";
defparam \Mux9~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~3 (
	.dataa(!ram_data_out2_13),
	.datab(!ram_data_out3_13),
	.datac(!ram_data_out0_13),
	.datad(!ram_data_out1_13),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~3 .extended_lut = "off";
defparam \Mux10~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux13~3 (
	.dataa(!ram_data_out2_10),
	.datab(!ram_data_out3_10),
	.datac(!ram_data_out0_10),
	.datad(!ram_data_out1_10),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~3 .extended_lut = "off";
defparam \Mux13~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux13~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux12~3 (
	.dataa(!ram_data_out2_11),
	.datab(!ram_data_out3_11),
	.datac(!ram_data_out0_11),
	.datad(!ram_data_out1_11),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux12~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~3 .extended_lut = "off";
defparam \Mux12~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux12~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~3 (
	.dataa(!ram_data_out2_12),
	.datab(!ram_data_out3_12),
	.datac(!ram_data_out0_12),
	.datad(!ram_data_out1_12),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~3 .extended_lut = "off";
defparam \Mux11~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux11~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!ram_data_out1_15),
	.datab(!ram_data_out2_15),
	.datac(!ram_data_out3_15),
	.datad(!ram_data_out0_15),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~1 (
	.dataa(!ram_data_out3_15),
	.datab(!ram_data_out0_15),
	.datac(!ram_data_out1_15),
	.datad(!ram_data_out2_15),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~1 .extended_lut = "off";
defparam \Mux8~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~2 (
	.dataa(!ram_data_out0_15),
	.datab(!ram_data_out1_15),
	.datac(!ram_data_out2_15),
	.datad(!ram_data_out3_15),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~2 .extended_lut = "off";
defparam \Mux8~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~3 (
	.dataa(!ram_data_out2_15),
	.datab(!ram_data_out3_15),
	.datac(!ram_data_out0_15),
	.datad(!ram_data_out1_15),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~3 .extended_lut = "off";
defparam \Mux8~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~0 (
	.dataa(!ram_data_out1_7),
	.datab(!ram_data_out2_7),
	.datac(!ram_data_out3_7),
	.datad(!ram_data_out0_7),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~0 .extended_lut = "off";
defparam \Mux40~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~0 (
	.dataa(!ram_data_out1_6),
	.datab(!ram_data_out2_6),
	.datac(!ram_data_out3_6),
	.datad(!ram_data_out0_6),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~0 .extended_lut = "off";
defparam \Mux41~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~0 (
	.dataa(!ram_data_out1_3),
	.datab(!ram_data_out2_3),
	.datac(!ram_data_out3_3),
	.datad(!ram_data_out0_3),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~0 .extended_lut = "off";
defparam \Mux44~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~0 (
	.dataa(!ram_data_out1_4),
	.datab(!ram_data_out2_4),
	.datac(!ram_data_out3_4),
	.datad(!ram_data_out0_4),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~0 .extended_lut = "off";
defparam \Mux43~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~0 (
	.dataa(!ram_data_out1_5),
	.datab(!ram_data_out2_5),
	.datac(!ram_data_out3_5),
	.datad(!ram_data_out0_5),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~0 .extended_lut = "off";
defparam \Mux42~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~1 (
	.dataa(!ram_data_out3_7),
	.datab(!ram_data_out0_7),
	.datac(!ram_data_out1_7),
	.datad(!ram_data_out2_7),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~1 .extended_lut = "off";
defparam \Mux40~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~1 (
	.dataa(!ram_data_out3_6),
	.datab(!ram_data_out0_6),
	.datac(!ram_data_out1_6),
	.datad(!ram_data_out2_6),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~1 .extended_lut = "off";
defparam \Mux41~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~1 (
	.dataa(!ram_data_out3_3),
	.datab(!ram_data_out0_3),
	.datac(!ram_data_out1_3),
	.datad(!ram_data_out2_3),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~1 .extended_lut = "off";
defparam \Mux44~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~1 (
	.dataa(!ram_data_out3_4),
	.datab(!ram_data_out0_4),
	.datac(!ram_data_out1_4),
	.datad(!ram_data_out2_4),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~1 .extended_lut = "off";
defparam \Mux43~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~1 (
	.dataa(!ram_data_out3_5),
	.datab(!ram_data_out0_5),
	.datac(!ram_data_out1_5),
	.datad(!ram_data_out2_5),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~1 .extended_lut = "off";
defparam \Mux42~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~2 (
	.dataa(!ram_data_out0_7),
	.datab(!ram_data_out1_7),
	.datac(!ram_data_out2_7),
	.datad(!ram_data_out3_7),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~2 .extended_lut = "off";
defparam \Mux40~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~2 (
	.dataa(!ram_data_out0_6),
	.datab(!ram_data_out1_6),
	.datac(!ram_data_out2_6),
	.datad(!ram_data_out3_6),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~2 .extended_lut = "off";
defparam \Mux41~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~2 (
	.dataa(!ram_data_out0_3),
	.datab(!ram_data_out1_3),
	.datac(!ram_data_out2_3),
	.datad(!ram_data_out3_3),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~2 .extended_lut = "off";
defparam \Mux44~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~2 (
	.dataa(!ram_data_out0_4),
	.datab(!ram_data_out1_4),
	.datac(!ram_data_out2_4),
	.datad(!ram_data_out3_4),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~2 .extended_lut = "off";
defparam \Mux43~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~2 (
	.dataa(!ram_data_out0_5),
	.datab(!ram_data_out1_5),
	.datac(!ram_data_out2_5),
	.datad(!ram_data_out3_5),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~2 .extended_lut = "off";
defparam \Mux42~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~3 (
	.dataa(!ram_data_out2_7),
	.datab(!ram_data_out3_7),
	.datac(!ram_data_out0_7),
	.datad(!ram_data_out1_7),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~3 .extended_lut = "off";
defparam \Mux40~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~3 (
	.dataa(!ram_data_out2_6),
	.datab(!ram_data_out3_6),
	.datac(!ram_data_out0_6),
	.datad(!ram_data_out1_6),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~3 .extended_lut = "off";
defparam \Mux41~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux44~3 (
	.dataa(!ram_data_out2_3),
	.datab(!ram_data_out3_3),
	.datac(!ram_data_out0_3),
	.datad(!ram_data_out1_3),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux44~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux44~3 .extended_lut = "off";
defparam \Mux44~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux44~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~3 (
	.dataa(!ram_data_out2_4),
	.datab(!ram_data_out3_4),
	.datac(!ram_data_out0_4),
	.datad(!ram_data_out1_4),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~3 .extended_lut = "off";
defparam \Mux43~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux43~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~3 (
	.dataa(!ram_data_out2_5),
	.datab(!ram_data_out3_5),
	.datac(!ram_data_out0_5),
	.datad(!ram_data_out1_5),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~3 .extended_lut = "off";
defparam \Mux42~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux42~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~0 (
	.dataa(!ram_data_out1_2),
	.datab(!ram_data_out2_2),
	.datac(!ram_data_out3_2),
	.datad(!ram_data_out0_2),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~0 .extended_lut = "off";
defparam \Mux45~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~1 (
	.dataa(!ram_data_out3_2),
	.datab(!ram_data_out0_2),
	.datac(!ram_data_out1_2),
	.datad(!ram_data_out2_2),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~1 .extended_lut = "off";
defparam \Mux45~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~2 (
	.dataa(!ram_data_out0_2),
	.datab(!ram_data_out1_2),
	.datac(!ram_data_out2_2),
	.datad(!ram_data_out3_2),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~2 .extended_lut = "off";
defparam \Mux45~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux45~3 (
	.dataa(!ram_data_out2_2),
	.datab(!ram_data_out3_2),
	.datac(!ram_data_out0_2),
	.datad(!ram_data_out1_2),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux45~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux45~3 .extended_lut = "off";
defparam \Mux45~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux45~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~0 (
	.dataa(!ram_data_out2_8),
	.datab(!ram_data_out3_8),
	.datac(!ram_data_out0_8),
	.datad(!ram_data_out1_8),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~0 .extended_lut = "off";
defparam \Mux15~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux15~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~0 (
	.dataa(!ram_data_out2_9),
	.datab(!ram_data_out3_9),
	.datac(!ram_data_out0_9),
	.datad(!ram_data_out1_9),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~0 .extended_lut = "off";
defparam \Mux14~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux14~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~1 (
	.dataa(!ram_data_out0_8),
	.datab(!ram_data_out1_8),
	.datac(!ram_data_out2_8),
	.datad(!ram_data_out3_8),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~1 .extended_lut = "off";
defparam \Mux15~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux15~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~1 (
	.dataa(!ram_data_out0_9),
	.datab(!ram_data_out1_9),
	.datac(!ram_data_out2_9),
	.datad(!ram_data_out3_9),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~1 .extended_lut = "off";
defparam \Mux14~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux14~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~0 (
	.dataa(!ram_data_out3_0),
	.datab(!ram_data_out0_0),
	.datac(!ram_data_out1_0),
	.datad(!ram_data_out2_0),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~0 .extended_lut = "off";
defparam \Mux47~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~0 (
	.dataa(!ram_data_out3_1),
	.datab(!ram_data_out0_1),
	.datac(!ram_data_out1_1),
	.datad(!ram_data_out2_1),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~0 .extended_lut = "off";
defparam \Mux46~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~1 (
	.dataa(!ram_data_out1_0),
	.datab(!ram_data_out2_0),
	.datac(!ram_data_out3_0),
	.datad(!ram_data_out0_0),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~1 .extended_lut = "off";
defparam \Mux47~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~1 (
	.dataa(!ram_data_out1_1),
	.datab(!ram_data_out2_1),
	.datac(!ram_data_out3_1),
	.datad(!ram_data_out0_1),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~1 .extended_lut = "off";
defparam \Mux46~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~2 (
	.dataa(!ram_data_out3_8),
	.datab(!ram_data_out0_8),
	.datac(!ram_data_out1_8),
	.datad(!ram_data_out2_8),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~2 .extended_lut = "off";
defparam \Mux15~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux15~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~2 (
	.dataa(!ram_data_out3_9),
	.datab(!ram_data_out0_9),
	.datac(!ram_data_out1_9),
	.datad(!ram_data_out2_9),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~2 .extended_lut = "off";
defparam \Mux14~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux14~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux15~3 (
	.dataa(!ram_data_out1_8),
	.datab(!ram_data_out2_8),
	.datac(!ram_data_out3_8),
	.datad(!ram_data_out0_8),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux15~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux15~3 .extended_lut = "off";
defparam \Mux15~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux15~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux14~3 (
	.dataa(!ram_data_out1_9),
	.datab(!ram_data_out2_9),
	.datac(!ram_data_out3_9),
	.datad(!ram_data_out0_9),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux14~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux14~3 .extended_lut = "off";
defparam \Mux14~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux14~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~2 (
	.dataa(!ram_data_out2_0),
	.datab(!ram_data_out3_0),
	.datac(!ram_data_out0_0),
	.datad(!ram_data_out1_0),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~2 .extended_lut = "off";
defparam \Mux47~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~2 (
	.dataa(!ram_data_out2_1),
	.datab(!ram_data_out3_1),
	.datac(!ram_data_out0_1),
	.datad(!ram_data_out1_1),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~2 .extended_lut = "off";
defparam \Mux46~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux47~3 (
	.dataa(!ram_data_out0_0),
	.datab(!ram_data_out1_0),
	.datac(!ram_data_out2_0),
	.datad(!ram_data_out3_0),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux47~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux47~3 .extended_lut = "off";
defparam \Mux47~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux47~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux46~3 (
	.dataa(!ram_data_out0_1),
	.datab(!ram_data_out1_1),
	.datac(!ram_data_out2_1),
	.datad(!ram_data_out3_1),
	.datae(!sw_r_tdl_0_4),
	.dataf(!sw_r_tdl_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux46~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux46~3 .extended_lut = "off";
defparam \Mux46~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux46~3 .shared_arith = "off";

endmodule

module IFFT_asj_fft_dataadgen (
	p_0,
	global_clock_enable,
	p_1,
	k_count_1,
	k_count_3,
	k_count_0,
	k_count_2,
	rd_addr_d_2,
	rd_addr_d_3,
	rd_addr_d_0,
	sw_0,
	rd_addr_c_0,
	rd_addr_b_1,
	sw_1,
	rd_addr_d_1,
	Mux1,
	Mux0,
	Mux11,
	Mux01,
	clk)/* synthesis synthesis_greybox=1 */;
input 	p_0;
input 	global_clock_enable;
input 	p_1;
input 	k_count_1;
input 	k_count_3;
input 	k_count_0;
input 	k_count_2;
output 	rd_addr_d_2;
output 	rd_addr_d_3;
output 	rd_addr_d_0;
output 	sw_0;
output 	rd_addr_c_0;
output 	rd_addr_b_1;
output 	sw_1;
output 	rd_addr_d_1;
output 	Mux1;
output 	Mux0;
output 	Mux11;
output 	Mux01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux4~0_combout ;
wire \Mux1~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;
wire \Mux0~0_combout ;
wire \Mux5~0_combout ;


dffeas \rd_addr_d[2] (
	.clk(clk),
	.d(k_count_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_d_2),
	.prn(vcc));
defparam \rd_addr_d[2] .is_wysiwyg = "true";
defparam \rd_addr_d[2] .power_up = "low";

dffeas \rd_addr_d[3] (
	.clk(clk),
	.d(k_count_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_d_3),
	.prn(vcc));
defparam \rd_addr_d[3] .is_wysiwyg = "true";
defparam \rd_addr_d[3] .power_up = "low";

dffeas \rd_addr_d[0] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_d_0),
	.prn(vcc));
defparam \rd_addr_d[0] .is_wysiwyg = "true";
defparam \rd_addr_d[0] .power_up = "low";

dffeas \sw[0] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(sw_0),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

dffeas \rd_addr_c[0] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_c_0),
	.prn(vcc));
defparam \rd_addr_c[0] .is_wysiwyg = "true";
defparam \rd_addr_c[0] .power_up = "low";

dffeas \rd_addr_b[1] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_b_1),
	.prn(vcc));
defparam \rd_addr_b[1] .is_wysiwyg = "true";
defparam \rd_addr_b[1] .power_up = "low";

dffeas \sw[1] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(sw_1),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

dffeas \rd_addr_d[1] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_d_1),
	.prn(vcc));
defparam \rd_addr_d[1] .is_wysiwyg = "true";
defparam \rd_addr_d[1] .power_up = "low";

cyclonev_lcell_comb \Mux1~1 (
	.dataa(!p_0),
	.datab(!k_count_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~1 .extended_lut = "off";
defparam \Mux1~1 .lut_mask = 64'h7777777777777777;
defparam \Mux1~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!p_0),
	.datab(!k_count_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'h7777777777777777;
defparam \Mux0~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~2 (
	.dataa(!p_0),
	.datab(!k_count_0),
	.datac(!k_count_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~2 .extended_lut = "off";
defparam \Mux1~2 .lut_mask = 64'h2727272727272727;
defparam \Mux1~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~2 (
	.dataa(!p_0),
	.datab(!k_count_1),
	.datac(!k_count_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~2 .extended_lut = "off";
defparam \Mux0~2 .lut_mask = 64'h2727272727272727;
defparam \Mux0~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!k_count_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!k_count_0),
	.datad(!k_count_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!k_count_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!k_count_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!k_count_1),
	.datad(!k_count_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!k_count_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Mux5~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_dft_bfp (
	next_block,
	reg_no_twiddle603,
	reg_no_twiddle607,
	reg_no_twiddle617,
	reg_no_twiddle613,
	reg_no_twiddle604,
	reg_no_twiddle614,
	reg_no_twiddle605,
	reg_no_twiddle615,
	reg_no_twiddle606,
	reg_no_twiddle616,
	reg_no_twiddle602,
	reg_no_twiddle612,
	reg_no_twiddle601,
	reg_no_twiddle611,
	tdl_arr_9,
	reg_no_twiddle600,
	reg_no_twiddle610,
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data007,
	twiddle_data107,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	twiddle_data207,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	global_clock_enable,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	lut_out_tmp_0,
	lut_out_tmp_1,
	lut_out_tmp_2,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_3_11,
	tdl_arr_7_11,
	tdl_arr_3_12,
	tdl_arr_7_12,
	tdl_arr_3_13,
	tdl_arr_7_13,
	tdl_arr_3_14,
	tdl_arr_7_14,
	tdl_arr_3_15,
	tdl_arr_7_15,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_4_12,
	tdl_arr_4_13,
	tdl_arr_4_14,
	tdl_arr_4_15,
	tdl_arr_5_1,
	tdl_arr_5_11,
	tdl_arr_5_12,
	tdl_arr_5_13,
	tdl_arr_5_14,
	tdl_arr_5_15,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_6_12,
	tdl_arr_6_13,
	tdl_arr_6_14,
	tdl_arr_6_15,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_2_12,
	tdl_arr_2_13,
	tdl_arr_2_14,
	tdl_arr_2_15,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_1_12,
	tdl_arr_1_13,
	tdl_arr_1_14,
	tdl_arr_1_15,
	tdl_arr_0_1,
	tdl_arr_0_11,
	tdl_arr_0_12,
	tdl_arr_0_13,
	tdl_arr_0_14,
	tdl_arr_0_15,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	ram_in_reg_6_1,
	ram_in_reg_5_1,
	ram_in_reg_2_1,
	ram_in_reg_3_1,
	ram_in_reg_4_1,
	ram_in_reg_6_3,
	ram_in_reg_5_3,
	ram_in_reg_2_3,
	ram_in_reg_3_3,
	ram_in_reg_4_3,
	ram_in_reg_6_0,
	ram_in_reg_5_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_6_2,
	ram_in_reg_5_2,
	ram_in_reg_2_2,
	ram_in_reg_3_2,
	ram_in_reg_4_2,
	ram_in_reg_7_1,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_2,
	ram_in_reg_7_5,
	ram_in_reg_6_5,
	ram_in_reg_3_5,
	ram_in_reg_4_5,
	ram_in_reg_5_5,
	ram_in_reg_7_7,
	ram_in_reg_6_7,
	ram_in_reg_3_7,
	ram_in_reg_4_7,
	ram_in_reg_5_7,
	ram_in_reg_7_4,
	ram_in_reg_6_4,
	ram_in_reg_3_4,
	ram_in_reg_4_4,
	ram_in_reg_5_4,
	ram_in_reg_7_6,
	ram_in_reg_6_6,
	ram_in_reg_3_6,
	ram_in_reg_4_6,
	ram_in_reg_5_6,
	ram_in_reg_2_5,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_6,
	ram_in_reg_0_2,
	ram_in_reg_1_2,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_0_7,
	ram_in_reg_1_7,
	ram_in_reg_0_5,
	ram_in_reg_1_5,
	ram_in_reg_0_3,
	ram_in_reg_1_3,
	ram_in_reg_0_1,
	ram_in_reg_1_1,
	ram_in_reg_0_6,
	ram_in_reg_1_6,
	ram_in_reg_0_4,
	ram_in_reg_1_4,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	next_block;
output 	reg_no_twiddle603;
output 	reg_no_twiddle607;
output 	reg_no_twiddle617;
output 	reg_no_twiddle613;
output 	reg_no_twiddle604;
output 	reg_no_twiddle614;
output 	reg_no_twiddle605;
output 	reg_no_twiddle615;
output 	reg_no_twiddle606;
output 	reg_no_twiddle616;
output 	reg_no_twiddle602;
output 	reg_no_twiddle612;
output 	reg_no_twiddle601;
output 	reg_no_twiddle611;
input 	tdl_arr_9;
output 	reg_no_twiddle600;
output 	reg_no_twiddle610;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data007;
input 	twiddle_data107;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	twiddle_data207;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	global_clock_enable;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
output 	lut_out_tmp_0;
output 	lut_out_tmp_1;
output 	lut_out_tmp_2;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_3_11;
output 	tdl_arr_7_11;
output 	tdl_arr_3_12;
output 	tdl_arr_7_12;
output 	tdl_arr_3_13;
output 	tdl_arr_7_13;
output 	tdl_arr_3_14;
output 	tdl_arr_7_14;
output 	tdl_arr_3_15;
output 	tdl_arr_7_15;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_4_12;
output 	tdl_arr_4_13;
output 	tdl_arr_4_14;
output 	tdl_arr_4_15;
output 	tdl_arr_5_1;
output 	tdl_arr_5_11;
output 	tdl_arr_5_12;
output 	tdl_arr_5_13;
output 	tdl_arr_5_14;
output 	tdl_arr_5_15;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_6_12;
output 	tdl_arr_6_13;
output 	tdl_arr_6_14;
output 	tdl_arr_6_15;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_2_12;
output 	tdl_arr_2_13;
output 	tdl_arr_2_14;
output 	tdl_arr_2_15;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_1_12;
output 	tdl_arr_1_13;
output 	tdl_arr_1_14;
output 	tdl_arr_1_15;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
output 	tdl_arr_0_12;
output 	tdl_arr_0_13;
output 	tdl_arr_0_14;
output 	tdl_arr_0_15;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	ram_in_reg_6_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_2_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_6_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_2_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_6_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_2_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_5;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_3_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_5_7;
input 	ram_in_reg_7_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_3_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_4;
input 	ram_in_reg_7_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_6;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_6;
input 	ram_in_reg_0_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_0_7;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_5;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_3;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_0_6;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_4;
input 	ram_in_reg_1_4;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \butterfly_st2[0][0][6]~q ;
wire \butterfly_st2[0][0][9]~q ;
wire \butterfly_st2[0][1][9]~q ;
wire \butterfly_st2[0][1][6]~q ;
wire \butterfly_st2[0][0][7]~q ;
wire \butterfly_st2[0][1][7]~q ;
wire \butterfly_st2[0][0][8]~q ;
wire \butterfly_st2[0][1][8]~q ;
wire \butterfly_st2[1][0][2]~q ;
wire \butterfly_st2[1][0][3]~q ;
wire \butterfly_st2[1][0][4]~q ;
wire \butterfly_st2[1][0][5]~q ;
wire \butterfly_st2[1][0][6]~q ;
wire \butterfly_st2[1][0][7]~q ;
wire \butterfly_st2[1][0][8]~q ;
wire \butterfly_st2[1][0][9]~q ;
wire \butterfly_st2[1][1][2]~q ;
wire \butterfly_st2[1][1][3]~q ;
wire \butterfly_st2[1][1][4]~q ;
wire \butterfly_st2[1][1][5]~q ;
wire \butterfly_st2[1][1][6]~q ;
wire \butterfly_st2[1][1][7]~q ;
wire \butterfly_st2[1][1][8]~q ;
wire \butterfly_st2[1][1][9]~q ;
wire \butterfly_st2[2][0][2]~q ;
wire \butterfly_st2[2][0][3]~q ;
wire \butterfly_st2[2][0][4]~q ;
wire \butterfly_st2[2][0][5]~q ;
wire \butterfly_st2[2][0][6]~q ;
wire \butterfly_st2[2][0][7]~q ;
wire \butterfly_st2[2][0][8]~q ;
wire \butterfly_st2[2][0][9]~q ;
wire \butterfly_st2[2][1][2]~q ;
wire \butterfly_st2[2][1][3]~q ;
wire \butterfly_st2[2][1][4]~q ;
wire \butterfly_st2[2][1][5]~q ;
wire \butterfly_st2[2][1][6]~q ;
wire \butterfly_st2[2][1][7]~q ;
wire \butterfly_st2[2][1][8]~q ;
wire \butterfly_st2[2][1][9]~q ;
wire \Add8~1_sumout ;
wire \Add8~2 ;
wire \butterfly_st2[0][0][5]~q ;
wire \Add8~5_sumout ;
wire \Add12~1_sumout ;
wire \Add12~5_sumout ;
wire \Add12~6 ;
wire \butterfly_st2[0][1][5]~q ;
wire \butterfly_st2[3][0][2]~q ;
wire \butterfly_st2[3][0][3]~q ;
wire \butterfly_st2[3][0][4]~q ;
wire \butterfly_st2[3][0][5]~q ;
wire \butterfly_st2[3][0][6]~q ;
wire \butterfly_st2[3][0][7]~q ;
wire \butterfly_st2[3][0][8]~q ;
wire \butterfly_st2[3][0][9]~q ;
wire \butterfly_st2[3][1][2]~q ;
wire \butterfly_st2[3][1][3]~q ;
wire \butterfly_st2[3][1][4]~q ;
wire \butterfly_st2[3][1][5]~q ;
wire \butterfly_st2[3][1][6]~q ;
wire \butterfly_st2[3][1][7]~q ;
wire \butterfly_st2[3][1][8]~q ;
wire \butterfly_st2[3][1][9]~q ;
wire \Add8~9_sumout ;
wire \Add8~10 ;
wire \Add12~9_sumout ;
wire \Add12~10 ;
wire \Add8~13_sumout ;
wire \Add8~14 ;
wire \Add12~13_sumout ;
wire \Add12~14 ;
wire \Add9~1_sumout ;
wire \Add9~2 ;
wire \butterfly_st2[1][0][1]~q ;
wire \Add9~5_sumout ;
wire \Add9~6 ;
wire \Add9~9_sumout ;
wire \Add9~10 ;
wire \Add9~13_sumout ;
wire \Add9~14 ;
wire \Add9~17_sumout ;
wire \Add9~18 ;
wire \Add9~21_sumout ;
wire \Add9~22 ;
wire \Add9~25_sumout ;
wire \Add9~26 ;
wire \Add9~29_sumout ;
wire \Add13~1_sumout ;
wire \Add13~2 ;
wire \Add13~3 ;
wire \butterfly_st2[1][1][1]~q ;
wire \Add13~5_sumout ;
wire \Add13~6 ;
wire \Add13~7 ;
wire \Add13~9_sumout ;
wire \Add13~10 ;
wire \Add13~11 ;
wire \Add13~13_sumout ;
wire \Add13~14 ;
wire \Add13~15 ;
wire \Add13~17_sumout ;
wire \Add13~18 ;
wire \Add13~19 ;
wire \Add13~21_sumout ;
wire \Add13~22 ;
wire \Add13~23 ;
wire \Add13~25_sumout ;
wire \Add13~26 ;
wire \Add13~27 ;
wire \Add13~29_sumout ;
wire \Add10~1_sumout ;
wire \Add10~2 ;
wire \Add10~3 ;
wire \butterfly_st2[2][0][1]~q ;
wire \Add10~5_sumout ;
wire \Add10~6 ;
wire \Add10~7 ;
wire \Add10~9_sumout ;
wire \Add10~10 ;
wire \Add10~11 ;
wire \Add10~13_sumout ;
wire \Add10~14 ;
wire \Add10~15 ;
wire \Add10~17_sumout ;
wire \Add10~18 ;
wire \Add10~19 ;
wire \Add10~21_sumout ;
wire \Add10~22 ;
wire \Add10~23 ;
wire \Add10~25_sumout ;
wire \Add10~26 ;
wire \Add10~27 ;
wire \Add10~29_sumout ;
wire \Add14~1_sumout ;
wire \Add14~2 ;
wire \Add14~3 ;
wire \butterfly_st2[2][1][1]~q ;
wire \Add14~5_sumout ;
wire \Add14~6 ;
wire \Add14~7 ;
wire \Add14~9_sumout ;
wire \Add14~10 ;
wire \Add14~11 ;
wire \Add14~13_sumout ;
wire \Add14~14 ;
wire \Add14~15 ;
wire \Add14~17_sumout ;
wire \Add14~18 ;
wire \Add14~19 ;
wire \Add14~21_sumout ;
wire \Add14~22 ;
wire \Add14~23 ;
wire \Add14~25_sumout ;
wire \Add14~26 ;
wire \Add14~27 ;
wire \Add14~29_sumout ;
wire \butterfly_st1[1][0][6]~q ;
wire \butterfly_st1[0][0][6]~q ;
wire \Add8~17_sumout ;
wire \Add8~18 ;
wire \butterfly_st2[0][0][4]~q ;
wire \butterfly_st1[1][0][8]~q ;
wire \butterfly_st1[0][0][8]~q ;
wire \butterfly_st1[1][1][8]~q ;
wire \butterfly_st1[0][1][8]~q ;
wire \butterfly_st1[1][1][6]~q ;
wire \butterfly_st1[0][1][6]~q ;
wire \Add12~17_sumout ;
wire \Add12~18 ;
wire \butterfly_st2[0][1][4]~q ;
wire \Add11~1_sumout ;
wire \Add11~2 ;
wire \Add11~3 ;
wire \butterfly_st2[3][0][1]~q ;
wire \Add11~5_sumout ;
wire \Add11~6 ;
wire \Add11~7 ;
wire \Add11~9_sumout ;
wire \Add11~10 ;
wire \Add11~11 ;
wire \Add11~13_sumout ;
wire \Add11~14 ;
wire \Add11~15 ;
wire \Add11~17_sumout ;
wire \Add11~18 ;
wire \Add11~19 ;
wire \Add11~21_sumout ;
wire \Add11~22 ;
wire \Add11~23 ;
wire \Add11~25_sumout ;
wire \Add11~26 ;
wire \Add11~27 ;
wire \Add11~29_sumout ;
wire \Add15~1_sumout ;
wire \Add15~2 ;
wire \butterfly_st2[3][1][1]~q ;
wire \Add15~5_sumout ;
wire \Add15~6 ;
wire \Add15~9_sumout ;
wire \Add15~10 ;
wire \Add15~13_sumout ;
wire \Add15~14 ;
wire \Add15~17_sumout ;
wire \Add15~18 ;
wire \Add15~21_sumout ;
wire \Add15~22 ;
wire \Add15~25_sumout ;
wire \Add15~26 ;
wire \Add15~29_sumout ;
wire \butterfly_st1[1][0][7]~q ;
wire \butterfly_st1[0][0][7]~q ;
wire \butterfly_st1[1][1][7]~q ;
wire \butterfly_st1[0][1][7]~q ;
wire \butterfly_st1[2][0][2]~q ;
wire \butterfly_st1[3][1][2]~q ;
wire \Add9~33_sumout ;
wire \Add9~34 ;
wire \butterfly_st2[1][0][0]~q ;
wire \butterfly_st1[2][0][3]~q ;
wire \butterfly_st1[3][1][3]~q ;
wire \butterfly_st1[2][0][4]~q ;
wire \butterfly_st1[3][1][4]~q ;
wire \butterfly_st1[2][0][5]~q ;
wire \butterfly_st1[3][1][5]~q ;
wire \butterfly_st1[2][0][6]~q ;
wire \butterfly_st1[3][1][6]~q ;
wire \butterfly_st1[2][0][7]~q ;
wire \butterfly_st1[3][1][7]~q ;
wire \butterfly_st1[2][0][8]~q ;
wire \butterfly_st1[3][1][8]~q ;
wire \butterfly_st1[3][0][2]~q ;
wire \butterfly_st1[2][1][2]~q ;
wire \Add13~33_sumout ;
wire \Add13~34 ;
wire \Add13~35 ;
wire \butterfly_st2[1][1][0]~q ;
wire \butterfly_st1[3][0][3]~q ;
wire \butterfly_st1[2][1][3]~q ;
wire \butterfly_st1[3][0][4]~q ;
wire \butterfly_st1[2][1][4]~q ;
wire \butterfly_st1[2][1][5]~q ;
wire \butterfly_st1[3][0][5]~q ;
wire \butterfly_st1[2][1][6]~q ;
wire \butterfly_st1[3][0][6]~q ;
wire \butterfly_st1[2][1][7]~q ;
wire \butterfly_st1[3][0][7]~q ;
wire \butterfly_st1[2][1][8]~q ;
wire \butterfly_st1[3][0][8]~q ;
wire \butterfly_st1[0][0][2]~q ;
wire \butterfly_st1[1][0][2]~q ;
wire \Add10~33_sumout ;
wire \Add10~34 ;
wire \Add10~35 ;
wire \butterfly_st2[2][0][0]~q ;
wire \butterfly_st1[0][0][3]~q ;
wire \butterfly_st1[1][0][3]~q ;
wire \butterfly_st1[0][0][4]~q ;
wire \butterfly_st1[1][0][4]~q ;
wire \butterfly_st1[0][0][5]~q ;
wire \butterfly_st1[1][0][5]~q ;
wire \butterfly_st1[0][1][2]~q ;
wire \butterfly_st1[1][1][2]~q ;
wire \Add14~33_sumout ;
wire \Add14~34 ;
wire \Add14~35 ;
wire \butterfly_st2[2][1][0]~q ;
wire \butterfly_st1[0][1][3]~q ;
wire \butterfly_st1[1][1][3]~q ;
wire \butterfly_st1[0][1][4]~q ;
wire \butterfly_st1[1][1][4]~q ;
wire \butterfly_st1[0][1][5]~q ;
wire \butterfly_st1[1][1][5]~q ;
wire \Add1~1_sumout ;
wire \Add1~2 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add8~21_sumout ;
wire \Add8~22 ;
wire \butterfly_st2[0][0][3]~q ;
wire \butterfly_st2[0][0][2]~q ;
wire \Add1~5_sumout ;
wire \Add0~5_sumout ;
wire \Add5~1_sumout ;
wire \Add4~1_sumout ;
wire \Add5~5_sumout ;
wire \Add5~6 ;
wire \Add4~5_sumout ;
wire \Add4~6 ;
wire \Add12~21_sumout ;
wire \Add12~22 ;
wire \butterfly_st2[0][1][3]~q ;
wire \butterfly_st2[0][1][2]~q ;
wire \Add11~33_sumout ;
wire \Add11~34 ;
wire \Add11~35 ;
wire \butterfly_st2[3][0][0]~q ;
wire \Add15~33_sumout ;
wire \Add15~34 ;
wire \butterfly_st2[3][1][0]~q ;
wire \Add1~9_sumout ;
wire \Add1~10 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add5~9_sumout ;
wire \Add5~10 ;
wire \Add4~9_sumout ;
wire \Add4~10 ;
wire \Add2~1_sumout ;
wire \Add2~2 ;
wire \Add2~3 ;
wire \Add7~1_sumout ;
wire \Add7~2 ;
wire \Add7~3 ;
wire \butterfly_st1[2][0][1]~q ;
wire \butterfly_st1[3][1][1]~q ;
wire \Add9~37_sumout ;
wire \Add9~38 ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add2~7 ;
wire \Add7~5_sumout ;
wire \Add7~6 ;
wire \Add7~7 ;
wire \Add2~9_sumout ;
wire \Add2~10 ;
wire \Add2~11 ;
wire \Add7~9_sumout ;
wire \Add7~10 ;
wire \Add7~11 ;
wire \Add2~13_sumout ;
wire \Add2~14 ;
wire \Add2~15 ;
wire \Add7~13_sumout ;
wire \Add7~14 ;
wire \Add7~15 ;
wire \Add2~17_sumout ;
wire \Add2~18 ;
wire \Add2~19 ;
wire \Add7~17_sumout ;
wire \Add7~18 ;
wire \Add7~19 ;
wire \Add2~21_sumout ;
wire \Add2~22 ;
wire \Add2~23 ;
wire \Add7~21_sumout ;
wire \Add7~22 ;
wire \Add7~23 ;
wire \Add2~25_sumout ;
wire \Add7~25_sumout ;
wire \Add3~1_sumout ;
wire \Add3~2 ;
wire \Add3~3 ;
wire \Add6~1_sumout ;
wire \Add6~2 ;
wire \Add6~3 ;
wire \butterfly_st1[3][0][1]~q ;
wire \butterfly_st1[2][1][1]~q ;
wire \Add13~37_sumout ;
wire \Add13~38 ;
wire \Add13~39 ;
wire \Add3~5_sumout ;
wire \Add3~6 ;
wire \Add3~7 ;
wire \Add6~5_sumout ;
wire \Add6~6 ;
wire \Add6~7 ;
wire \Add3~9_sumout ;
wire \Add3~10 ;
wire \Add3~11 ;
wire \Add6~9_sumout ;
wire \Add6~10 ;
wire \Add6~11 ;
wire \Add6~13_sumout ;
wire \Add6~14 ;
wire \Add6~15 ;
wire \Add3~13_sumout ;
wire \Add3~14 ;
wire \Add3~15 ;
wire \Add6~17_sumout ;
wire \Add6~18 ;
wire \Add6~19 ;
wire \Add3~17_sumout ;
wire \Add3~18 ;
wire \Add3~19 ;
wire \Add6~21_sumout ;
wire \Add6~22 ;
wire \Add6~23 ;
wire \Add3~21_sumout ;
wire \Add3~22 ;
wire \Add3~23 ;
wire \Add6~25_sumout ;
wire \Add3~25_sumout ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add1~13_sumout ;
wire \Add1~14 ;
wire \butterfly_st1[0][0][1]~q ;
wire \butterfly_st1[1][0][1]~q ;
wire \Add10~37_sumout ;
wire \Add10~38 ;
wire \Add10~39 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add1~17_sumout ;
wire \Add1~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add1~21_sumout ;
wire \Add1~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add1~25_sumout ;
wire \Add1~26 ;
wire \Add4~13_sumout ;
wire \Add4~14 ;
wire \Add5~13_sumout ;
wire \Add5~14 ;
wire \butterfly_st1[0][1][1]~q ;
wire \butterfly_st1[1][1][1]~q ;
wire \Add14~37_sumout ;
wire \Add14~38 ;
wire \Add14~39 ;
wire \Add4~17_sumout ;
wire \Add4~18 ;
wire \Add5~17_sumout ;
wire \Add5~18 ;
wire \Add4~21_sumout ;
wire \Add4~22 ;
wire \Add5~21_sumout ;
wire \Add5~22 ;
wire \Add4~25_sumout ;
wire \Add4~26 ;
wire \Add5~25_sumout ;
wire \Add5~26 ;
wire \Add8~25_sumout ;
wire \Add8~26 ;
wire \Add8~29_sumout ;
wire \Add8~30 ;
wire \butterfly_st2[0][0][1]~q ;
wire \Add12~25_sumout ;
wire \Add12~26 ;
wire \Add12~29_sumout ;
wire \Add12~30 ;
wire \butterfly_st2[0][1][1]~q ;
wire \Add11~37_sumout ;
wire \Add11~38 ;
wire \Add11~39 ;
wire \Add15~37_sumout ;
wire \Add15~38 ;
wire \gen_disc:bfp_scale|r_array_out[2][2]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][2]~q ;
wire \Add2~29_sumout ;
wire \Add2~30 ;
wire \Add2~31 ;
wire \gen_disc:bfp_scale|i_array_out[3][2]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][2]~q ;
wire \Add7~29_sumout ;
wire \Add7~30 ;
wire \Add7~31 ;
wire \butterfly_st1[2][0][0]~q ;
wire \butterfly_st1[3][1][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][2]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][2]~q ;
wire \Add3~29_sumout ;
wire \Add3~30 ;
wire \Add3~31 ;
wire \gen_disc:bfp_scale|i_array_out[2][2]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][2]~q ;
wire \Add6~29_sumout ;
wire \Add6~30 ;
wire \Add6~31 ;
wire \butterfly_st1[3][0][0]~q ;
wire \butterfly_st1[2][1][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][3]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][3]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][4]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][4]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][5]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][5]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][5]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add1~29_sumout ;
wire \Add1~30 ;
wire \butterfly_st1[0][0][0]~q ;
wire \butterfly_st1[1][0][0]~q ;
wire \Add4~29_sumout ;
wire \Add4~30 ;
wire \Add5~29_sumout ;
wire \Add5~30 ;
wire \butterfly_st1[0][1][0]~q ;
wire \butterfly_st1[1][1][0]~q ;
wire \Add8~33_sumout ;
wire \Add8~34 ;
wire \butterfly_st2[0][0][0]~q ;
wire \Add12~33_sumout ;
wire \Add12~34 ;
wire \butterfly_st2[0][1][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][1]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][1]~q ;
wire \Add2~33_sumout ;
wire \Add2~34 ;
wire \Add2~35 ;
wire \gen_disc:bfp_scale|i_array_out[3][1]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][1]~q ;
wire \Add7~33_sumout ;
wire \Add7~34 ;
wire \Add7~35 ;
wire \gen_disc:bfp_scale|r_array_out[3][1]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][1]~q ;
wire \Add3~33_sumout ;
wire \Add3~34 ;
wire \Add3~35 ;
wire \gen_disc:bfp_scale|i_array_out[2][1]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][1]~q ;
wire \Add6~33_sumout ;
wire \Add6~34 ;
wire \Add6~35 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add1~33_sumout ;
wire \Add1~34 ;
wire \Add4~33_sumout ;
wire \Add4~34 ;
wire \Add5~33_sumout ;
wire \Add5~34 ;
wire \Add8~37_sumout ;
wire \Add8~38 ;
wire \Add12~37_sumout ;
wire \Add12~38 ;
wire \gen_disc:bfp_scale|r_array_out[2][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][0]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][0]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][0]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][6]~q ;
wire \gen_disc:bfp_scale|r_array_out[1][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[3][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[0][7]~q ;
wire \gen_disc:bfp_scale|r_array_out[2][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][7]~q ;
wire \gen_disc:bfp_scale|i_array_out[1][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[3][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[0][6]~q ;
wire \gen_disc:bfp_scale|i_array_out[2][6]~q ;
wire \Add16~30 ;
wire \Add16~26 ;
wire \Add16~22 ;
wire \Add16~1_sumout ;
wire \reg_no_twiddle[0][0][3]~q ;
wire \reg_no_twiddle[1][0][3]~q ;
wire \reg_no_twiddle[2][0][3]~q ;
wire \reg_no_twiddle[3][0][3]~q ;
wire \reg_no_twiddle[4][0][3]~q ;
wire \reg_no_twiddle[5][0][3]~q ;
wire \Add16~2 ;
wire \Add16~10 ;
wire \Add16~14 ;
wire \Add16~18 ;
wire \Add16~5_sumout ;
wire \reg_no_twiddle[0][0][7]~q ;
wire \reg_no_twiddle[1][0][7]~q ;
wire \reg_no_twiddle[2][0][7]~q ;
wire \reg_no_twiddle[3][0][7]~q ;
wire \reg_no_twiddle[4][0][7]~q ;
wire \reg_no_twiddle[5][0][7]~q ;
wire \Add17~30 ;
wire \Add17~26 ;
wire \Add17~22 ;
wire \Add17~6 ;
wire \Add17~10 ;
wire \Add17~14 ;
wire \Add17~18 ;
wire \Add17~1_sumout ;
wire \reg_no_twiddle[0][1][7]~q ;
wire \reg_no_twiddle[1][1][7]~q ;
wire \reg_no_twiddle[2][1][7]~q ;
wire \reg_no_twiddle[3][1][7]~q ;
wire \reg_no_twiddle[4][1][7]~q ;
wire \reg_no_twiddle[5][1][7]~q ;
wire \Add17~5_sumout ;
wire \reg_no_twiddle[0][1][3]~q ;
wire \reg_no_twiddle[1][1][3]~q ;
wire \reg_no_twiddle[2][1][3]~q ;
wire \reg_no_twiddle[3][1][3]~q ;
wire \reg_no_twiddle[4][1][3]~q ;
wire \reg_no_twiddle[5][1][3]~q ;
wire \Add16~9_sumout ;
wire \reg_no_twiddle[0][0][4]~q ;
wire \reg_no_twiddle[1][0][4]~q ;
wire \reg_no_twiddle[2][0][4]~q ;
wire \reg_no_twiddle[3][0][4]~q ;
wire \reg_no_twiddle[4][0][4]~q ;
wire \reg_no_twiddle[5][0][4]~q ;
wire \Add17~9_sumout ;
wire \reg_no_twiddle[0][1][4]~q ;
wire \reg_no_twiddle[1][1][4]~q ;
wire \reg_no_twiddle[2][1][4]~q ;
wire \reg_no_twiddle[3][1][4]~q ;
wire \reg_no_twiddle[4][1][4]~q ;
wire \reg_no_twiddle[5][1][4]~q ;
wire \Add16~13_sumout ;
wire \reg_no_twiddle[0][0][5]~q ;
wire \reg_no_twiddle[1][0][5]~q ;
wire \reg_no_twiddle[2][0][5]~q ;
wire \reg_no_twiddle[3][0][5]~q ;
wire \reg_no_twiddle[4][0][5]~q ;
wire \reg_no_twiddle[5][0][5]~q ;
wire \Add17~13_sumout ;
wire \reg_no_twiddle[0][1][5]~q ;
wire \reg_no_twiddle[1][1][5]~q ;
wire \reg_no_twiddle[2][1][5]~q ;
wire \reg_no_twiddle[3][1][5]~q ;
wire \reg_no_twiddle[4][1][5]~q ;
wire \reg_no_twiddle[5][1][5]~q ;
wire \Add16~17_sumout ;
wire \reg_no_twiddle[0][0][6]~q ;
wire \reg_no_twiddle[1][0][6]~q ;
wire \reg_no_twiddle[2][0][6]~q ;
wire \reg_no_twiddle[3][0][6]~q ;
wire \reg_no_twiddle[4][0][6]~q ;
wire \reg_no_twiddle[5][0][6]~q ;
wire \Add17~17_sumout ;
wire \reg_no_twiddle[0][1][6]~q ;
wire \reg_no_twiddle[1][1][6]~q ;
wire \reg_no_twiddle[2][1][6]~q ;
wire \reg_no_twiddle[3][1][6]~q ;
wire \reg_no_twiddle[4][1][6]~q ;
wire \reg_no_twiddle[5][1][6]~q ;
wire \Add16~21_sumout ;
wire \reg_no_twiddle[0][0][2]~q ;
wire \reg_no_twiddle[1][0][2]~q ;
wire \reg_no_twiddle[2][0][2]~q ;
wire \reg_no_twiddle[3][0][2]~q ;
wire \reg_no_twiddle[4][0][2]~q ;
wire \reg_no_twiddle[5][0][2]~q ;
wire \Add17~21_sumout ;
wire \reg_no_twiddle[0][1][2]~q ;
wire \reg_no_twiddle[1][1][2]~q ;
wire \reg_no_twiddle[2][1][2]~q ;
wire \reg_no_twiddle[3][1][2]~q ;
wire \reg_no_twiddle[4][1][2]~q ;
wire \reg_no_twiddle[5][1][2]~q ;
wire \Add16~25_sumout ;
wire \reg_no_twiddle[0][0][1]~q ;
wire \reg_no_twiddle[1][0][1]~q ;
wire \reg_no_twiddle[2][0][1]~q ;
wire \reg_no_twiddle[3][0][1]~q ;
wire \reg_no_twiddle[4][0][1]~q ;
wire \reg_no_twiddle[5][0][1]~q ;
wire \Add17~25_sumout ;
wire \reg_no_twiddle[0][1][1]~q ;
wire \reg_no_twiddle[1][1][1]~q ;
wire \reg_no_twiddle[2][1][1]~q ;
wire \reg_no_twiddle[3][1][1]~q ;
wire \reg_no_twiddle[4][1][1]~q ;
wire \reg_no_twiddle[5][1][1]~q ;
wire \Add16~29_sumout ;
wire \reg_no_twiddle[0][0][0]~q ;
wire \reg_no_twiddle[1][0][0]~q ;
wire \reg_no_twiddle[2][0][0]~q ;
wire \reg_no_twiddle[3][0][0]~q ;
wire \reg_no_twiddle[4][0][0]~q ;
wire \reg_no_twiddle[5][0][0]~q ;
wire \Add17~29_sumout ;
wire \reg_no_twiddle[0][1][0]~q ;
wire \reg_no_twiddle[1][1][0]~q ;
wire \reg_no_twiddle[2][1][0]~q ;
wire \reg_no_twiddle[3][1][0]~q ;
wire \reg_no_twiddle[4][1][0]~q ;
wire \reg_no_twiddle[5][1][0]~q ;


IFFT_apn_fft_cmult_cpx2 \gen_da2:cm1 (
	.twiddle_data010(twiddle_data010),
	.twiddle_data011(twiddle_data011),
	.twiddle_data012(twiddle_data012),
	.twiddle_data013(twiddle_data013),
	.twiddle_data014(twiddle_data014),
	.twiddle_data015(twiddle_data015),
	.twiddle_data016(twiddle_data016),
	.twiddle_data017(twiddle_data017),
	.twiddle_data007(twiddle_data007),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_3_11(tdl_arr_3_13),
	.tdl_arr_7_11(tdl_arr_7_13),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_4_11(tdl_arr_4_13),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_5_11(tdl_arr_5_13),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_6_11(tdl_arr_6_13),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_2_11(tdl_arr_2_14),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_1_11(tdl_arr_1_14),
	.tdl_arr_0_1(tdl_arr_0_11),
	.tdl_arr_0_11(tdl_arr_0_14),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.twiddle_data000(twiddle_data000),
	.twiddle_data001(twiddle_data001),
	.twiddle_data002(twiddle_data002),
	.twiddle_data003(twiddle_data003),
	.twiddle_data004(twiddle_data004),
	.twiddle_data005(twiddle_data005),
	.twiddle_data006(twiddle_data006),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk),
	.reset(reset_n));

IFFT_asj_fft_bfp_i \gen_disc:bfp_scale (
	.r_array_out_2_2(\gen_disc:bfp_scale|r_array_out[2][2]~q ),
	.r_array_out_2_0(\gen_disc:bfp_scale|r_array_out[0][2]~q ),
	.i_array_out_2_3(\gen_disc:bfp_scale|i_array_out[3][2]~q ),
	.i_array_out_2_1(\gen_disc:bfp_scale|i_array_out[1][2]~q ),
	.r_array_out_3_0(\gen_disc:bfp_scale|r_array_out[0][3]~q ),
	.r_array_out_3_2(\gen_disc:bfp_scale|r_array_out[2][3]~q ),
	.i_array_out_3_1(\gen_disc:bfp_scale|i_array_out[1][3]~q ),
	.i_array_out_3_3(\gen_disc:bfp_scale|i_array_out[3][3]~q ),
	.r_array_out_4_2(\gen_disc:bfp_scale|r_array_out[2][4]~q ),
	.r_array_out_4_0(\gen_disc:bfp_scale|r_array_out[0][4]~q ),
	.i_array_out_4_3(\gen_disc:bfp_scale|i_array_out[3][4]~q ),
	.i_array_out_4_1(\gen_disc:bfp_scale|i_array_out[1][4]~q ),
	.r_array_out_5_2(\gen_disc:bfp_scale|r_array_out[2][5]~q ),
	.r_array_out_5_0(\gen_disc:bfp_scale|r_array_out[0][5]~q ),
	.i_array_out_5_3(\gen_disc:bfp_scale|i_array_out[3][5]~q ),
	.i_array_out_5_1(\gen_disc:bfp_scale|i_array_out[1][5]~q ),
	.r_array_out_2_3(\gen_disc:bfp_scale|r_array_out[3][2]~q ),
	.r_array_out_2_1(\gen_disc:bfp_scale|r_array_out[1][2]~q ),
	.i_array_out_2_2(\gen_disc:bfp_scale|i_array_out[2][2]~q ),
	.i_array_out_2_0(\gen_disc:bfp_scale|i_array_out[0][2]~q ),
	.r_array_out_3_3(\gen_disc:bfp_scale|r_array_out[3][3]~q ),
	.r_array_out_3_1(\gen_disc:bfp_scale|r_array_out[1][3]~q ),
	.i_array_out_3_0(\gen_disc:bfp_scale|i_array_out[0][3]~q ),
	.i_array_out_3_2(\gen_disc:bfp_scale|i_array_out[2][3]~q ),
	.r_array_out_4_3(\gen_disc:bfp_scale|r_array_out[3][4]~q ),
	.r_array_out_4_1(\gen_disc:bfp_scale|r_array_out[1][4]~q ),
	.i_array_out_4_2(\gen_disc:bfp_scale|i_array_out[2][4]~q ),
	.i_array_out_4_0(\gen_disc:bfp_scale|i_array_out[0][4]~q ),
	.i_array_out_5_2(\gen_disc:bfp_scale|i_array_out[2][5]~q ),
	.i_array_out_5_0(\gen_disc:bfp_scale|i_array_out[0][5]~q ),
	.r_array_out_5_3(\gen_disc:bfp_scale|r_array_out[3][5]~q ),
	.r_array_out_5_1(\gen_disc:bfp_scale|r_array_out[1][5]~q ),
	.r_array_out_1_0(\gen_disc:bfp_scale|r_array_out[0][1]~q ),
	.r_array_out_1_2(\gen_disc:bfp_scale|r_array_out[2][1]~q ),
	.i_array_out_1_3(\gen_disc:bfp_scale|i_array_out[3][1]~q ),
	.i_array_out_1_1(\gen_disc:bfp_scale|i_array_out[1][1]~q ),
	.r_array_out_1_3(\gen_disc:bfp_scale|r_array_out[3][1]~q ),
	.r_array_out_1_1(\gen_disc:bfp_scale|r_array_out[1][1]~q ),
	.i_array_out_1_2(\gen_disc:bfp_scale|i_array_out[2][1]~q ),
	.i_array_out_1_0(\gen_disc:bfp_scale|i_array_out[0][1]~q ),
	.r_array_out_0_2(\gen_disc:bfp_scale|r_array_out[2][0]~q ),
	.r_array_out_0_0(\gen_disc:bfp_scale|r_array_out[0][0]~q ),
	.i_array_out_0_1(\gen_disc:bfp_scale|i_array_out[1][0]~q ),
	.i_array_out_0_3(\gen_disc:bfp_scale|i_array_out[3][0]~q ),
	.r_array_out_0_3(\gen_disc:bfp_scale|r_array_out[3][0]~q ),
	.r_array_out_0_1(\gen_disc:bfp_scale|r_array_out[1][0]~q ),
	.i_array_out_0_2(\gen_disc:bfp_scale|i_array_out[2][0]~q ),
	.i_array_out_0_0(\gen_disc:bfp_scale|i_array_out[0][0]~q ),
	.global_clock_enable(global_clock_enable),
	.slb_last_0(slb_last_0),
	.slb_last_1(slb_last_1),
	.slb_last_2(slb_last_2),
	.r_array_out_6_1(\gen_disc:bfp_scale|r_array_out[1][6]~q ),
	.r_array_out_6_3(\gen_disc:bfp_scale|r_array_out[3][6]~q ),
	.r_array_out_6_0(\gen_disc:bfp_scale|r_array_out[0][6]~q ),
	.r_array_out_6_2(\gen_disc:bfp_scale|r_array_out[2][6]~q ),
	.r_array_out_7_1(\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.r_array_out_7_3(\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.r_array_out_7_0(\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.r_array_out_7_2(\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.i_array_out_7_1(\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.i_array_out_7_3(\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.i_array_out_7_0(\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.i_array_out_7_2(\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.i_array_out_6_1(\gen_disc:bfp_scale|i_array_out[1][6]~q ),
	.i_array_out_6_3(\gen_disc:bfp_scale|i_array_out[3][6]~q ),
	.i_array_out_6_0(\gen_disc:bfp_scale|i_array_out[0][6]~q ),
	.i_array_out_6_2(\gen_disc:bfp_scale|i_array_out[2][6]~q ),
	.ram_in_reg_6_1(ram_in_reg_6_1),
	.ram_in_reg_5_1(ram_in_reg_5_1),
	.ram_in_reg_2_1(ram_in_reg_2_1),
	.ram_in_reg_3_1(ram_in_reg_3_1),
	.ram_in_reg_4_1(ram_in_reg_4_1),
	.ram_in_reg_6_3(ram_in_reg_6_3),
	.ram_in_reg_5_3(ram_in_reg_5_3),
	.ram_in_reg_2_3(ram_in_reg_2_3),
	.ram_in_reg_3_3(ram_in_reg_3_3),
	.ram_in_reg_4_3(ram_in_reg_4_3),
	.ram_in_reg_6_0(ram_in_reg_6_0),
	.ram_in_reg_5_0(ram_in_reg_5_0),
	.ram_in_reg_2_0(ram_in_reg_2_0),
	.ram_in_reg_3_0(ram_in_reg_3_0),
	.ram_in_reg_4_0(ram_in_reg_4_0),
	.ram_in_reg_6_2(ram_in_reg_6_2),
	.ram_in_reg_5_2(ram_in_reg_5_2),
	.ram_in_reg_2_2(ram_in_reg_2_2),
	.ram_in_reg_3_2(ram_in_reg_3_2),
	.ram_in_reg_4_2(ram_in_reg_4_2),
	.ram_in_reg_7_1(ram_in_reg_7_1),
	.ram_in_reg_7_3(ram_in_reg_7_3),
	.ram_in_reg_7_0(ram_in_reg_7_0),
	.ram_in_reg_7_2(ram_in_reg_7_2),
	.ram_in_reg_7_5(ram_in_reg_7_5),
	.ram_in_reg_6_5(ram_in_reg_6_5),
	.ram_in_reg_3_5(ram_in_reg_3_5),
	.ram_in_reg_4_5(ram_in_reg_4_5),
	.ram_in_reg_5_5(ram_in_reg_5_5),
	.ram_in_reg_7_7(ram_in_reg_7_7),
	.ram_in_reg_6_7(ram_in_reg_6_7),
	.ram_in_reg_3_7(ram_in_reg_3_7),
	.ram_in_reg_4_7(ram_in_reg_4_7),
	.ram_in_reg_5_7(ram_in_reg_5_7),
	.ram_in_reg_7_4(ram_in_reg_7_4),
	.ram_in_reg_6_4(ram_in_reg_6_4),
	.ram_in_reg_3_4(ram_in_reg_3_4),
	.ram_in_reg_4_4(ram_in_reg_4_4),
	.ram_in_reg_5_4(ram_in_reg_5_4),
	.ram_in_reg_7_6(ram_in_reg_7_6),
	.ram_in_reg_6_6(ram_in_reg_6_6),
	.ram_in_reg_3_6(ram_in_reg_3_6),
	.ram_in_reg_4_6(ram_in_reg_4_6),
	.ram_in_reg_5_6(ram_in_reg_5_6),
	.ram_in_reg_2_5(ram_in_reg_2_5),
	.ram_in_reg_2_7(ram_in_reg_2_7),
	.ram_in_reg_2_4(ram_in_reg_2_4),
	.ram_in_reg_2_6(ram_in_reg_2_6),
	.ram_in_reg_0_2(ram_in_reg_0_2),
	.ram_in_reg_1_2(ram_in_reg_1_2),
	.ram_in_reg_0_0(ram_in_reg_0_0),
	.ram_in_reg_1_0(ram_in_reg_1_0),
	.ram_in_reg_0_7(ram_in_reg_0_7),
	.ram_in_reg_1_7(ram_in_reg_1_7),
	.ram_in_reg_0_5(ram_in_reg_0_5),
	.ram_in_reg_1_5(ram_in_reg_1_5),
	.ram_in_reg_0_3(ram_in_reg_0_3),
	.ram_in_reg_1_3(ram_in_reg_1_3),
	.ram_in_reg_0_1(ram_in_reg_0_1),
	.ram_in_reg_1_1(ram_in_reg_1_1),
	.ram_in_reg_0_6(ram_in_reg_0_6),
	.ram_in_reg_1_6(ram_in_reg_1_6),
	.ram_in_reg_0_4(ram_in_reg_0_4),
	.ram_in_reg_1_4(ram_in_reg_1_4),
	.clk(clk));

IFFT_asj_fft_bfp_o \gen_disc:bfp_detect (
	.next_block(next_block),
	.reg_no_twiddle603(reg_no_twiddle603),
	.reg_no_twiddle607(reg_no_twiddle607),
	.reg_no_twiddle617(reg_no_twiddle617),
	.reg_no_twiddle613(reg_no_twiddle613),
	.reg_no_twiddle604(reg_no_twiddle604),
	.reg_no_twiddle614(reg_no_twiddle614),
	.reg_no_twiddle605(reg_no_twiddle605),
	.reg_no_twiddle615(reg_no_twiddle615),
	.reg_no_twiddle606(reg_no_twiddle606),
	.reg_no_twiddle616(reg_no_twiddle616),
	.tdl_arr_9(tdl_arr_9),
	.global_clock_enable(global_clock_enable),
	.lut_out_tmp_0(lut_out_tmp_0),
	.lut_out_tmp_1(lut_out_tmp_1),
	.lut_out_tmp_2(lut_out_tmp_2),
	.tdl_arr_3_1(tdl_arr_3_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_3_11(tdl_arr_3_11),
	.tdl_arr_7_11(tdl_arr_7_11),
	.tdl_arr_3_12(tdl_arr_3_12),
	.tdl_arr_7_12(tdl_arr_7_12),
	.tdl_arr_3_13(tdl_arr_3_13),
	.tdl_arr_7_13(tdl_arr_7_13),
	.tdl_arr_3_14(tdl_arr_3_14),
	.tdl_arr_7_14(tdl_arr_7_14),
	.tdl_arr_3_15(tdl_arr_3_15),
	.tdl_arr_7_15(tdl_arr_7_15),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_4_11(tdl_arr_4_11),
	.tdl_arr_4_12(tdl_arr_4_12),
	.tdl_arr_4_13(tdl_arr_4_13),
	.tdl_arr_4_14(tdl_arr_4_14),
	.tdl_arr_4_15(tdl_arr_4_15),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_5_11(tdl_arr_5_11),
	.tdl_arr_5_12(tdl_arr_5_12),
	.tdl_arr_5_13(tdl_arr_5_13),
	.tdl_arr_5_14(tdl_arr_5_14),
	.tdl_arr_5_15(tdl_arr_5_15),
	.tdl_arr_6_1(tdl_arr_6_1),
	.tdl_arr_6_11(tdl_arr_6_11),
	.tdl_arr_6_12(tdl_arr_6_12),
	.tdl_arr_6_13(tdl_arr_6_13),
	.tdl_arr_6_14(tdl_arr_6_14),
	.tdl_arr_6_15(tdl_arr_6_15),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_pround_13 \gen_full_rnd:gen_rounding_blk:3:u1 (
	.butterfly_st2312(\butterfly_st2[3][1][2]~q ),
	.butterfly_st2313(\butterfly_st2[3][1][3]~q ),
	.butterfly_st2314(\butterfly_st2[3][1][4]~q ),
	.butterfly_st2315(\butterfly_st2[3][1][5]~q ),
	.butterfly_st2316(\butterfly_st2[3][1][6]~q ),
	.butterfly_st2317(\butterfly_st2[3][1][7]~q ),
	.butterfly_st2318(\butterfly_st2[3][1][8]~q ),
	.butterfly_st2319(\butterfly_st2[3][1][9]~q ),
	.butterfly_st2311(\butterfly_st2[3][1][1]~q ),
	.butterfly_st2310(\butterfly_st2[3][1][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk));

IFFT_asj_fft_pround_12 \gen_full_rnd:gen_rounding_blk:3:u0 (
	.butterfly_st2302(\butterfly_st2[3][0][2]~q ),
	.butterfly_st2303(\butterfly_st2[3][0][3]~q ),
	.butterfly_st2304(\butterfly_st2[3][0][4]~q ),
	.butterfly_st2305(\butterfly_st2[3][0][5]~q ),
	.butterfly_st2306(\butterfly_st2[3][0][6]~q ),
	.butterfly_st2307(\butterfly_st2[3][0][7]~q ),
	.butterfly_st2308(\butterfly_st2[3][0][8]~q ),
	.butterfly_st2309(\butterfly_st2[3][0][9]~q ),
	.butterfly_st2301(\butterfly_st2[3][0][1]~q ),
	.butterfly_st2300(\butterfly_st2[3][0][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk));

IFFT_asj_fft_pround_11 \gen_full_rnd:gen_rounding_blk:2:u1 (
	.butterfly_st2212(\butterfly_st2[2][1][2]~q ),
	.butterfly_st2213(\butterfly_st2[2][1][3]~q ),
	.butterfly_st2214(\butterfly_st2[2][1][4]~q ),
	.butterfly_st2215(\butterfly_st2[2][1][5]~q ),
	.butterfly_st2216(\butterfly_st2[2][1][6]~q ),
	.butterfly_st2217(\butterfly_st2[2][1][7]~q ),
	.butterfly_st2218(\butterfly_st2[2][1][8]~q ),
	.butterfly_st2219(\butterfly_st2[2][1][9]~q ),
	.butterfly_st2211(\butterfly_st2[2][1][1]~q ),
	.butterfly_st2210(\butterfly_st2[2][1][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk));

IFFT_asj_fft_pround_10 \gen_full_rnd:gen_rounding_blk:2:u0 (
	.butterfly_st2202(\butterfly_st2[2][0][2]~q ),
	.butterfly_st2203(\butterfly_st2[2][0][3]~q ),
	.butterfly_st2204(\butterfly_st2[2][0][4]~q ),
	.butterfly_st2205(\butterfly_st2[2][0][5]~q ),
	.butterfly_st2206(\butterfly_st2[2][0][6]~q ),
	.butterfly_st2207(\butterfly_st2[2][0][7]~q ),
	.butterfly_st2208(\butterfly_st2[2][0][8]~q ),
	.butterfly_st2209(\butterfly_st2[2][0][9]~q ),
	.butterfly_st2201(\butterfly_st2[2][0][1]~q ),
	.butterfly_st2200(\butterfly_st2[2][0][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk));

IFFT_asj_fft_pround_9 \gen_full_rnd:gen_rounding_blk:1:u1 (
	.butterfly_st2112(\butterfly_st2[1][1][2]~q ),
	.butterfly_st2113(\butterfly_st2[1][1][3]~q ),
	.butterfly_st2114(\butterfly_st2[1][1][4]~q ),
	.butterfly_st2115(\butterfly_st2[1][1][5]~q ),
	.butterfly_st2116(\butterfly_st2[1][1][6]~q ),
	.butterfly_st2117(\butterfly_st2[1][1][7]~q ),
	.butterfly_st2118(\butterfly_st2[1][1][8]~q ),
	.butterfly_st2119(\butterfly_st2[1][1][9]~q ),
	.butterfly_st2111(\butterfly_st2[1][1][1]~q ),
	.butterfly_st2110(\butterfly_st2[1][1][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk));

IFFT_asj_fft_pround_8 \gen_full_rnd:gen_rounding_blk:1:u0 (
	.butterfly_st2102(\butterfly_st2[1][0][2]~q ),
	.butterfly_st2103(\butterfly_st2[1][0][3]~q ),
	.butterfly_st2104(\butterfly_st2[1][0][4]~q ),
	.butterfly_st2105(\butterfly_st2[1][0][5]~q ),
	.butterfly_st2106(\butterfly_st2[1][0][6]~q ),
	.butterfly_st2107(\butterfly_st2[1][0][7]~q ),
	.butterfly_st2108(\butterfly_st2[1][0][8]~q ),
	.butterfly_st2109(\butterfly_st2[1][0][9]~q ),
	.butterfly_st2101(\butterfly_st2[1][0][1]~q ),
	.butterfly_st2100(\butterfly_st2[1][0][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk));

IFFT_asj_fft_pround_7 \gen_full_rnd:gen_rounding_blk:0:u1 (
	.butterfly_st2019(\butterfly_st2[0][1][9]~q ),
	.butterfly_st2016(\butterfly_st2[0][1][6]~q ),
	.butterfly_st2017(\butterfly_st2[0][1][7]~q ),
	.butterfly_st2018(\butterfly_st2[0][1][8]~q ),
	.butterfly_st2015(\butterfly_st2[0][1][5]~q ),
	.butterfly_st2014(\butterfly_st2[0][1][4]~q ),
	.butterfly_st2013(\butterfly_st2[0][1][3]~q ),
	.butterfly_st2012(\butterfly_st2[0][1][2]~q ),
	.butterfly_st2011(\butterfly_st2[0][1][1]~q ),
	.butterfly_st2010(\butterfly_st2[0][1][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.clk(clk));

IFFT_asj_fft_pround_6 \gen_full_rnd:gen_rounding_blk:0:u0 (
	.butterfly_st2006(\butterfly_st2[0][0][6]~q ),
	.butterfly_st2009(\butterfly_st2[0][0][9]~q ),
	.butterfly_st2007(\butterfly_st2[0][0][7]~q ),
	.butterfly_st2008(\butterfly_st2[0][0][8]~q ),
	.butterfly_st2005(\butterfly_st2[0][0][5]~q ),
	.butterfly_st2004(\butterfly_st2[0][0][4]~q ),
	.butterfly_st2003(\butterfly_st2[0][0][3]~q ),
	.butterfly_st2002(\butterfly_st2[0][0][2]~q ),
	.butterfly_st2001(\butterfly_st2[0][0][1]~q ),
	.butterfly_st2000(\butterfly_st2[0][0][0]~q ),
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.clk(clk));

IFFT_apn_fft_cmult_cpx2_2 \gen_da2:cm3 (
	.twiddle_data207(twiddle_data207),
	.twiddle_data210(twiddle_data210),
	.twiddle_data211(twiddle_data211),
	.twiddle_data212(twiddle_data212),
	.twiddle_data213(twiddle_data213),
	.twiddle_data214(twiddle_data214),
	.twiddle_data215(twiddle_data215),
	.twiddle_data216(twiddle_data216),
	.twiddle_data217(twiddle_data217),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_14),
	.tdl_arr_7_1(tdl_arr_7_14),
	.tdl_arr_3_11(tdl_arr_3_15),
	.tdl_arr_7_11(tdl_arr_7_15),
	.tdl_arr_4_1(tdl_arr_4_14),
	.tdl_arr_4_11(tdl_arr_4_15),
	.tdl_arr_5_1(tdl_arr_5_14),
	.tdl_arr_5_11(tdl_arr_5_15),
	.tdl_arr_6_1(tdl_arr_6_14),
	.tdl_arr_6_11(tdl_arr_6_15),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_2_11(tdl_arr_2_13),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_1_11(tdl_arr_1_13),
	.tdl_arr_0_1(tdl_arr_0_1),
	.tdl_arr_0_11(tdl_arr_0_13),
	.twiddle_data200(twiddle_data200),
	.twiddle_data201(twiddle_data201),
	.twiddle_data202(twiddle_data202),
	.twiddle_data203(twiddle_data203),
	.twiddle_data204(twiddle_data204),
	.twiddle_data205(twiddle_data205),
	.twiddle_data206(twiddle_data206),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk),
	.reset(reset_n));

IFFT_apn_fft_cmult_cpx2_1 \gen_da2:cm2 (
	.twiddle_data107(twiddle_data107),
	.twiddle_data110(twiddle_data110),
	.twiddle_data111(twiddle_data111),
	.twiddle_data112(twiddle_data112),
	.twiddle_data113(twiddle_data113),
	.twiddle_data114(twiddle_data114),
	.twiddle_data115(twiddle_data115),
	.twiddle_data116(twiddle_data116),
	.twiddle_data117(twiddle_data117),
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_3_11(tdl_arr_3_12),
	.tdl_arr_7_11(tdl_arr_7_12),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_4_11(tdl_arr_4_12),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_5_11(tdl_arr_5_12),
	.tdl_arr_6_1(tdl_arr_6_11),
	.tdl_arr_6_11(tdl_arr_6_12),
	.tdl_arr_2_1(tdl_arr_2_12),
	.tdl_arr_2_11(tdl_arr_2_15),
	.tdl_arr_1_1(tdl_arr_1_12),
	.tdl_arr_1_11(tdl_arr_1_15),
	.tdl_arr_0_1(tdl_arr_0_12),
	.tdl_arr_0_11(tdl_arr_0_15),
	.twiddle_data100(twiddle_data100),
	.twiddle_data101(twiddle_data101),
	.twiddle_data102(twiddle_data102),
	.twiddle_data103(twiddle_data103),
	.twiddle_data104(twiddle_data104),
	.twiddle_data105(twiddle_data105),
	.twiddle_data106(twiddle_data106),
	.pipeline_dffe_2(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_21(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk),
	.reset(reset_n));

dffeas \butterfly_st2[0][0][6] (
	.clk(clk),
	.d(\Add8~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][6] .power_up = "low";

dffeas \butterfly_st2[0][0][9] (
	.clk(clk),
	.d(\Add8~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][9] .power_up = "low";

dffeas \butterfly_st2[0][1][9] (
	.clk(clk),
	.d(\Add12~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][9] .power_up = "low";

dffeas \butterfly_st2[0][1][6] (
	.clk(clk),
	.d(\Add12~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][6] .power_up = "low";

dffeas \butterfly_st2[0][0][7] (
	.clk(clk),
	.d(\Add8~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][7] .power_up = "low";

dffeas \butterfly_st2[0][1][7] (
	.clk(clk),
	.d(\Add12~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][7] .power_up = "low";

dffeas \butterfly_st2[0][0][8] (
	.clk(clk),
	.d(\Add8~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][8] .power_up = "low";

dffeas \butterfly_st2[0][1][8] (
	.clk(clk),
	.d(\Add12~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][8] .power_up = "low";

dffeas \butterfly_st2[1][0][2] (
	.clk(clk),
	.d(\Add9~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][2] .power_up = "low";

dffeas \butterfly_st2[1][0][3] (
	.clk(clk),
	.d(\Add9~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][3] .power_up = "low";

dffeas \butterfly_st2[1][0][4] (
	.clk(clk),
	.d(\Add9~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][4] .power_up = "low";

dffeas \butterfly_st2[1][0][5] (
	.clk(clk),
	.d(\Add9~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][5] .power_up = "low";

dffeas \butterfly_st2[1][0][6] (
	.clk(clk),
	.d(\Add9~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][6] .power_up = "low";

dffeas \butterfly_st2[1][0][7] (
	.clk(clk),
	.d(\Add9~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][7] .power_up = "low";

dffeas \butterfly_st2[1][0][8] (
	.clk(clk),
	.d(\Add9~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][8] .power_up = "low";

dffeas \butterfly_st2[1][0][9] (
	.clk(clk),
	.d(\Add9~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][9] .power_up = "low";

dffeas \butterfly_st2[1][1][2] (
	.clk(clk),
	.d(\Add13~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][2] .power_up = "low";

dffeas \butterfly_st2[1][1][3] (
	.clk(clk),
	.d(\Add13~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][3] .power_up = "low";

dffeas \butterfly_st2[1][1][4] (
	.clk(clk),
	.d(\Add13~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][4] .power_up = "low";

dffeas \butterfly_st2[1][1][5] (
	.clk(clk),
	.d(\Add13~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][5] .power_up = "low";

dffeas \butterfly_st2[1][1][6] (
	.clk(clk),
	.d(\Add13~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][6] .power_up = "low";

dffeas \butterfly_st2[1][1][7] (
	.clk(clk),
	.d(\Add13~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][7] .power_up = "low";

dffeas \butterfly_st2[1][1][8] (
	.clk(clk),
	.d(\Add13~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][8] .power_up = "low";

dffeas \butterfly_st2[1][1][9] (
	.clk(clk),
	.d(\Add13~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][9] .power_up = "low";

dffeas \butterfly_st2[2][0][2] (
	.clk(clk),
	.d(\Add10~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][2] .power_up = "low";

dffeas \butterfly_st2[2][0][3] (
	.clk(clk),
	.d(\Add10~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][3] .power_up = "low";

dffeas \butterfly_st2[2][0][4] (
	.clk(clk),
	.d(\Add10~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][4] .power_up = "low";

dffeas \butterfly_st2[2][0][5] (
	.clk(clk),
	.d(\Add10~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][5] .power_up = "low";

dffeas \butterfly_st2[2][0][6] (
	.clk(clk),
	.d(\Add10~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][6] .power_up = "low";

dffeas \butterfly_st2[2][0][7] (
	.clk(clk),
	.d(\Add10~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][7] .power_up = "low";

dffeas \butterfly_st2[2][0][8] (
	.clk(clk),
	.d(\Add10~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][8] .power_up = "low";

dffeas \butterfly_st2[2][0][9] (
	.clk(clk),
	.d(\Add10~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][9] .power_up = "low";

dffeas \butterfly_st2[2][1][2] (
	.clk(clk),
	.d(\Add14~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][2] .power_up = "low";

dffeas \butterfly_st2[2][1][3] (
	.clk(clk),
	.d(\Add14~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][3] .power_up = "low";

dffeas \butterfly_st2[2][1][4] (
	.clk(clk),
	.d(\Add14~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][4] .power_up = "low";

dffeas \butterfly_st2[2][1][5] (
	.clk(clk),
	.d(\Add14~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][5] .power_up = "low";

dffeas \butterfly_st2[2][1][6] (
	.clk(clk),
	.d(\Add14~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][6] .power_up = "low";

dffeas \butterfly_st2[2][1][7] (
	.clk(clk),
	.d(\Add14~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][7] .power_up = "low";

dffeas \butterfly_st2[2][1][8] (
	.clk(clk),
	.d(\Add14~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][8] .power_up = "low";

dffeas \butterfly_st2[2][1][9] (
	.clk(clk),
	.d(\Add14~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][9] .power_up = "low";

cyclonev_lcell_comb \Add8~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][6]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][6]~q ),
	.datag(gnd),
	.cin(\Add8~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~1_sumout ),
	.cout(\Add8~2 ),
	.shareout());
defparam \Add8~1 .extended_lut = "off";
defparam \Add8~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~1 .shared_arith = "off";

dffeas \butterfly_st2[0][0][5] (
	.clk(clk),
	.d(\Add8~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][5] .power_up = "low";

cyclonev_lcell_comb \Add8~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][8]~q ),
	.datag(gnd),
	.cin(\Add8~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~5_sumout ),
	.cout(),
	.shareout());
defparam \Add8~5 .extended_lut = "off";
defparam \Add8~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~5 .shared_arith = "off";

cyclonev_lcell_comb \Add12~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][8]~q ),
	.datag(gnd),
	.cin(\Add12~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~1_sumout ),
	.cout(),
	.shareout());
defparam \Add12~1 .extended_lut = "off";
defparam \Add12~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~1 .shared_arith = "off";

cyclonev_lcell_comb \Add12~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][6]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][6]~q ),
	.datag(gnd),
	.cin(\Add12~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~5_sumout ),
	.cout(\Add12~6 ),
	.shareout());
defparam \Add12~5 .extended_lut = "off";
defparam \Add12~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~5 .shared_arith = "off";

dffeas \butterfly_st2[0][1][5] (
	.clk(clk),
	.d(\Add12~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][5] .power_up = "low";

dffeas \butterfly_st2[3][0][2] (
	.clk(clk),
	.d(\Add11~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][2] .power_up = "low";

dffeas \butterfly_st2[3][0][3] (
	.clk(clk),
	.d(\Add11~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][3] .power_up = "low";

dffeas \butterfly_st2[3][0][4] (
	.clk(clk),
	.d(\Add11~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][4] .power_up = "low";

dffeas \butterfly_st2[3][0][5] (
	.clk(clk),
	.d(\Add11~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][5] .power_up = "low";

dffeas \butterfly_st2[3][0][6] (
	.clk(clk),
	.d(\Add11~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][6] .power_up = "low";

dffeas \butterfly_st2[3][0][7] (
	.clk(clk),
	.d(\Add11~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][7] .power_up = "low";

dffeas \butterfly_st2[3][0][8] (
	.clk(clk),
	.d(\Add11~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][8] .power_up = "low";

dffeas \butterfly_st2[3][0][9] (
	.clk(clk),
	.d(\Add11~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][9] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][9] .power_up = "low";

dffeas \butterfly_st2[3][1][2] (
	.clk(clk),
	.d(\Add15~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][2] .power_up = "low";

dffeas \butterfly_st2[3][1][3] (
	.clk(clk),
	.d(\Add15~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][3] .power_up = "low";

dffeas \butterfly_st2[3][1][4] (
	.clk(clk),
	.d(\Add15~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][4] .power_up = "low";

dffeas \butterfly_st2[3][1][5] (
	.clk(clk),
	.d(\Add15~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][5] .power_up = "low";

dffeas \butterfly_st2[3][1][6] (
	.clk(clk),
	.d(\Add15~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][6] .power_up = "low";

dffeas \butterfly_st2[3][1][7] (
	.clk(clk),
	.d(\Add15~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][7] .power_up = "low";

dffeas \butterfly_st2[3][1][8] (
	.clk(clk),
	.d(\Add15~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][8] .power_up = "low";

dffeas \butterfly_st2[3][1][9] (
	.clk(clk),
	.d(\Add15~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][9]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][9] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][9] .power_up = "low";

cyclonev_lcell_comb \Add8~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][7]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][7]~q ),
	.datag(gnd),
	.cin(\Add8~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~9_sumout ),
	.cout(\Add8~10 ),
	.shareout());
defparam \Add8~9 .extended_lut = "off";
defparam \Add8~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~9 .shared_arith = "off";

cyclonev_lcell_comb \Add12~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][7]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][7]~q ),
	.datag(gnd),
	.cin(\Add12~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~9_sumout ),
	.cout(\Add12~10 ),
	.shareout());
defparam \Add12~9 .extended_lut = "off";
defparam \Add12~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~9 .shared_arith = "off";

cyclonev_lcell_comb \Add8~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][8]~q ),
	.datag(gnd),
	.cin(\Add8~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~13_sumout ),
	.cout(\Add8~14 ),
	.shareout());
defparam \Add8~13 .extended_lut = "off";
defparam \Add8~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~13 .shared_arith = "off";

cyclonev_lcell_comb \Add12~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][8]~q ),
	.datag(gnd),
	.cin(\Add12~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~13_sumout ),
	.cout(\Add12~14 ),
	.shareout());
defparam \Add12~13 .extended_lut = "off";
defparam \Add12~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~13 .shared_arith = "off";

cyclonev_lcell_comb \Add9~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][2]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][2]~q ),
	.datag(gnd),
	.cin(\Add9~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~1_sumout ),
	.cout(\Add9~2 ),
	.shareout());
defparam \Add9~1 .extended_lut = "off";
defparam \Add9~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~1 .shared_arith = "off";

dffeas \butterfly_st2[1][0][1] (
	.clk(clk),
	.d(\Add9~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][1] .power_up = "low";

cyclonev_lcell_comb \Add9~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][3]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][3]~q ),
	.datag(gnd),
	.cin(\Add9~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~5_sumout ),
	.cout(\Add9~6 ),
	.shareout());
defparam \Add9~5 .extended_lut = "off";
defparam \Add9~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~5 .shared_arith = "off";

cyclonev_lcell_comb \Add9~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][4]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][4]~q ),
	.datag(gnd),
	.cin(\Add9~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~9_sumout ),
	.cout(\Add9~10 ),
	.shareout());
defparam \Add9~9 .extended_lut = "off";
defparam \Add9~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~9 .shared_arith = "off";

cyclonev_lcell_comb \Add9~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][5]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][5]~q ),
	.datag(gnd),
	.cin(\Add9~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~13_sumout ),
	.cout(\Add9~14 ),
	.shareout());
defparam \Add9~13 .extended_lut = "off";
defparam \Add9~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~13 .shared_arith = "off";

cyclonev_lcell_comb \Add9~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][6]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][6]~q ),
	.datag(gnd),
	.cin(\Add9~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~17_sumout ),
	.cout(\Add9~18 ),
	.shareout());
defparam \Add9~17 .extended_lut = "off";
defparam \Add9~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~17 .shared_arith = "off";

cyclonev_lcell_comb \Add9~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][7]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][7]~q ),
	.datag(gnd),
	.cin(\Add9~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~21_sumout ),
	.cout(\Add9~22 ),
	.shareout());
defparam \Add9~21 .extended_lut = "off";
defparam \Add9~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~21 .shared_arith = "off";

cyclonev_lcell_comb \Add9~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][8]~q ),
	.datag(gnd),
	.cin(\Add9~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~25_sumout ),
	.cout(\Add9~26 ),
	.shareout());
defparam \Add9~25 .extended_lut = "off";
defparam \Add9~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~25 .shared_arith = "off";

cyclonev_lcell_comb \Add9~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][8]~q ),
	.datag(gnd),
	.cin(\Add9~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~29_sumout ),
	.cout(),
	.shareout());
defparam \Add9~29 .extended_lut = "off";
defparam \Add9~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~29 .shared_arith = "off";

cyclonev_lcell_comb \Add13~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][0][2]~q ),
	.datad(!\butterfly_st1[2][1][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~34 ),
	.sharein(\Add13~35 ),
	.combout(),
	.sumout(\Add13~1_sumout ),
	.cout(\Add13~2 ),
	.shareout(\Add13~3 ));
defparam \Add13~1 .extended_lut = "off";
defparam \Add13~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add13~1 .shared_arith = "on";

dffeas \butterfly_st2[1][1][1] (
	.clk(clk),
	.d(\Add13~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][1] .power_up = "low";

cyclonev_lcell_comb \Add13~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][0][3]~q ),
	.datad(!\butterfly_st1[2][1][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~2 ),
	.sharein(\Add13~3 ),
	.combout(),
	.sumout(\Add13~5_sumout ),
	.cout(\Add13~6 ),
	.shareout(\Add13~7 ));
defparam \Add13~5 .extended_lut = "off";
defparam \Add13~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add13~5 .shared_arith = "on";

cyclonev_lcell_comb \Add13~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][0][4]~q ),
	.datad(!\butterfly_st1[2][1][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~6 ),
	.sharein(\Add13~7 ),
	.combout(),
	.sumout(\Add13~9_sumout ),
	.cout(\Add13~10 ),
	.shareout(\Add13~11 ));
defparam \Add13~9 .extended_lut = "off";
defparam \Add13~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add13~9 .shared_arith = "on";

cyclonev_lcell_comb \Add13~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[2][1][5]~q ),
	.datad(!\butterfly_st1[3][0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~10 ),
	.sharein(\Add13~11 ),
	.combout(),
	.sumout(\Add13~13_sumout ),
	.cout(\Add13~14 ),
	.shareout(\Add13~15 ));
defparam \Add13~13 .extended_lut = "off";
defparam \Add13~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add13~13 .shared_arith = "on";

cyclonev_lcell_comb \Add13~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[2][1][6]~q ),
	.datad(!\butterfly_st1[3][0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~14 ),
	.sharein(\Add13~15 ),
	.combout(),
	.sumout(\Add13~17_sumout ),
	.cout(\Add13~18 ),
	.shareout(\Add13~19 ));
defparam \Add13~17 .extended_lut = "off";
defparam \Add13~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add13~17 .shared_arith = "on";

cyclonev_lcell_comb \Add13~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[2][1][7]~q ),
	.datad(!\butterfly_st1[3][0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~18 ),
	.sharein(\Add13~19 ),
	.combout(),
	.sumout(\Add13~21_sumout ),
	.cout(\Add13~22 ),
	.shareout(\Add13~23 ));
defparam \Add13~21 .extended_lut = "off";
defparam \Add13~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add13~21 .shared_arith = "on";

cyclonev_lcell_comb \Add13~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[2][1][8]~q ),
	.datad(!\butterfly_st1[3][0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~22 ),
	.sharein(\Add13~23 ),
	.combout(),
	.sumout(\Add13~25_sumout ),
	.cout(\Add13~26 ),
	.shareout(\Add13~27 ));
defparam \Add13~25 .extended_lut = "off";
defparam \Add13~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add13~25 .shared_arith = "on";

cyclonev_lcell_comb \Add13~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[2][1][8]~q ),
	.datad(!\butterfly_st1[3][0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~26 ),
	.sharein(\Add13~27 ),
	.combout(),
	.sumout(\Add13~29_sumout ),
	.cout(),
	.shareout());
defparam \Add13~29 .extended_lut = "off";
defparam \Add13~29 .lut_mask = 64'h0000000000000FF0;
defparam \Add13~29 .shared_arith = "on";

cyclonev_lcell_comb \Add10~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][2]~q ),
	.datad(!\butterfly_st1[1][0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~34 ),
	.sharein(\Add10~35 ),
	.combout(),
	.sumout(\Add10~1_sumout ),
	.cout(\Add10~2 ),
	.shareout(\Add10~3 ));
defparam \Add10~1 .extended_lut = "off";
defparam \Add10~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~1 .shared_arith = "on";

dffeas \butterfly_st2[2][0][1] (
	.clk(clk),
	.d(\Add10~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][1] .power_up = "low";

cyclonev_lcell_comb \Add10~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][3]~q ),
	.datad(!\butterfly_st1[1][0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~2 ),
	.sharein(\Add10~3 ),
	.combout(),
	.sumout(\Add10~5_sumout ),
	.cout(\Add10~6 ),
	.shareout(\Add10~7 ));
defparam \Add10~5 .extended_lut = "off";
defparam \Add10~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~5 .shared_arith = "on";

cyclonev_lcell_comb \Add10~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][4]~q ),
	.datad(!\butterfly_st1[1][0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~6 ),
	.sharein(\Add10~7 ),
	.combout(),
	.sumout(\Add10~9_sumout ),
	.cout(\Add10~10 ),
	.shareout(\Add10~11 ));
defparam \Add10~9 .extended_lut = "off";
defparam \Add10~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~9 .shared_arith = "on";

cyclonev_lcell_comb \Add10~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][5]~q ),
	.datad(!\butterfly_st1[1][0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~10 ),
	.sharein(\Add10~11 ),
	.combout(),
	.sumout(\Add10~13_sumout ),
	.cout(\Add10~14 ),
	.shareout(\Add10~15 ));
defparam \Add10~13 .extended_lut = "off";
defparam \Add10~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~13 .shared_arith = "on";

cyclonev_lcell_comb \Add10~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][6]~q ),
	.datad(!\butterfly_st1[1][0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~14 ),
	.sharein(\Add10~15 ),
	.combout(),
	.sumout(\Add10~17_sumout ),
	.cout(\Add10~18 ),
	.shareout(\Add10~19 ));
defparam \Add10~17 .extended_lut = "off";
defparam \Add10~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~17 .shared_arith = "on";

cyclonev_lcell_comb \Add10~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][7]~q ),
	.datad(!\butterfly_st1[1][0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~18 ),
	.sharein(\Add10~19 ),
	.combout(),
	.sumout(\Add10~21_sumout ),
	.cout(\Add10~22 ),
	.shareout(\Add10~23 ));
defparam \Add10~21 .extended_lut = "off";
defparam \Add10~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~21 .shared_arith = "on";

cyclonev_lcell_comb \Add10~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][8]~q ),
	.datad(!\butterfly_st1[1][0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~22 ),
	.sharein(\Add10~23 ),
	.combout(),
	.sumout(\Add10~25_sumout ),
	.cout(\Add10~26 ),
	.shareout(\Add10~27 ));
defparam \Add10~25 .extended_lut = "off";
defparam \Add10~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~25 .shared_arith = "on";

cyclonev_lcell_comb \Add10~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][8]~q ),
	.datad(!\butterfly_st1[1][0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~26 ),
	.sharein(\Add10~27 ),
	.combout(),
	.sumout(\Add10~29_sumout ),
	.cout(),
	.shareout());
defparam \Add10~29 .extended_lut = "off";
defparam \Add10~29 .lut_mask = 64'h0000000000000FF0;
defparam \Add10~29 .shared_arith = "on";

cyclonev_lcell_comb \Add14~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][2]~q ),
	.datad(!\butterfly_st1[1][1][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~34 ),
	.sharein(\Add14~35 ),
	.combout(),
	.sumout(\Add14~1_sumout ),
	.cout(\Add14~2 ),
	.shareout(\Add14~3 ));
defparam \Add14~1 .extended_lut = "off";
defparam \Add14~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~1 .shared_arith = "on";

dffeas \butterfly_st2[2][1][1] (
	.clk(clk),
	.d(\Add14~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][1] .power_up = "low";

cyclonev_lcell_comb \Add14~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][3]~q ),
	.datad(!\butterfly_st1[1][1][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~2 ),
	.sharein(\Add14~3 ),
	.combout(),
	.sumout(\Add14~5_sumout ),
	.cout(\Add14~6 ),
	.shareout(\Add14~7 ));
defparam \Add14~5 .extended_lut = "off";
defparam \Add14~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~5 .shared_arith = "on";

cyclonev_lcell_comb \Add14~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][4]~q ),
	.datad(!\butterfly_st1[1][1][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~6 ),
	.sharein(\Add14~7 ),
	.combout(),
	.sumout(\Add14~9_sumout ),
	.cout(\Add14~10 ),
	.shareout(\Add14~11 ));
defparam \Add14~9 .extended_lut = "off";
defparam \Add14~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~9 .shared_arith = "on";

cyclonev_lcell_comb \Add14~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][5]~q ),
	.datad(!\butterfly_st1[1][1][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~10 ),
	.sharein(\Add14~11 ),
	.combout(),
	.sumout(\Add14~13_sumout ),
	.cout(\Add14~14 ),
	.shareout(\Add14~15 ));
defparam \Add14~13 .extended_lut = "off";
defparam \Add14~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~13 .shared_arith = "on";

cyclonev_lcell_comb \Add14~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][6]~q ),
	.datad(!\butterfly_st1[1][1][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~14 ),
	.sharein(\Add14~15 ),
	.combout(),
	.sumout(\Add14~17_sumout ),
	.cout(\Add14~18 ),
	.shareout(\Add14~19 ));
defparam \Add14~17 .extended_lut = "off";
defparam \Add14~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~17 .shared_arith = "on";

cyclonev_lcell_comb \Add14~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][7]~q ),
	.datad(!\butterfly_st1[1][1][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~18 ),
	.sharein(\Add14~19 ),
	.combout(),
	.sumout(\Add14~21_sumout ),
	.cout(\Add14~22 ),
	.shareout(\Add14~23 ));
defparam \Add14~21 .extended_lut = "off";
defparam \Add14~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~21 .shared_arith = "on";

cyclonev_lcell_comb \Add14~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][8]~q ),
	.datad(!\butterfly_st1[1][1][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~22 ),
	.sharein(\Add14~23 ),
	.combout(),
	.sumout(\Add14~25_sumout ),
	.cout(\Add14~26 ),
	.shareout(\Add14~27 ));
defparam \Add14~25 .extended_lut = "off";
defparam \Add14~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~25 .shared_arith = "on";

cyclonev_lcell_comb \Add14~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][8]~q ),
	.datad(!\butterfly_st1[1][1][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~26 ),
	.sharein(\Add14~27 ),
	.combout(),
	.sumout(\Add14~29_sumout ),
	.cout(),
	.shareout());
defparam \Add14~29 .extended_lut = "off";
defparam \Add14~29 .lut_mask = 64'h0000000000000FF0;
defparam \Add14~29 .shared_arith = "on";

dffeas \butterfly_st1[1][0][6] (
	.clk(clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][6] .power_up = "low";

dffeas \butterfly_st1[0][0][6] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][6] .power_up = "low";

cyclonev_lcell_comb \Add8~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][5]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][5]~q ),
	.datag(gnd),
	.cin(\Add8~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~17_sumout ),
	.cout(\Add8~18 ),
	.shareout());
defparam \Add8~17 .extended_lut = "off";
defparam \Add8~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~17 .shared_arith = "off";

dffeas \butterfly_st2[0][0][4] (
	.clk(clk),
	.d(\Add8~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][4] .power_up = "low";

dffeas \butterfly_st1[1][0][8] (
	.clk(clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][8] .power_up = "low";

dffeas \butterfly_st1[0][0][8] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][8] .power_up = "low";

dffeas \butterfly_st1[1][1][8] (
	.clk(clk),
	.d(\Add5~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][8] .power_up = "low";

dffeas \butterfly_st1[0][1][8] (
	.clk(clk),
	.d(\Add4~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][8] .power_up = "low";

dffeas \butterfly_st1[1][1][6] (
	.clk(clk),
	.d(\Add5~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][6] .power_up = "low";

dffeas \butterfly_st1[0][1][6] (
	.clk(clk),
	.d(\Add4~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][6] .power_up = "low";

cyclonev_lcell_comb \Add12~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][5]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][5]~q ),
	.datag(gnd),
	.cin(\Add12~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~17_sumout ),
	.cout(\Add12~18 ),
	.shareout());
defparam \Add12~17 .extended_lut = "off";
defparam \Add12~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~17 .shared_arith = "off";

dffeas \butterfly_st2[0][1][4] (
	.clk(clk),
	.d(\Add12~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][4] .power_up = "low";

cyclonev_lcell_comb \Add11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][2]~q ),
	.datad(!\butterfly_st1[2][0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~34 ),
	.sharein(\Add11~35 ),
	.combout(),
	.sumout(\Add11~1_sumout ),
	.cout(\Add11~2 ),
	.shareout(\Add11~3 ));
defparam \Add11~1 .extended_lut = "off";
defparam \Add11~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~1 .shared_arith = "on";

dffeas \butterfly_st2[3][0][1] (
	.clk(clk),
	.d(\Add11~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][1] .power_up = "low";

cyclonev_lcell_comb \Add11~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][3]~q ),
	.datad(!\butterfly_st1[2][0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~2 ),
	.sharein(\Add11~3 ),
	.combout(),
	.sumout(\Add11~5_sumout ),
	.cout(\Add11~6 ),
	.shareout(\Add11~7 ));
defparam \Add11~5 .extended_lut = "off";
defparam \Add11~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~5 .shared_arith = "on";

cyclonev_lcell_comb \Add11~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][4]~q ),
	.datad(!\butterfly_st1[2][0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~6 ),
	.sharein(\Add11~7 ),
	.combout(),
	.sumout(\Add11~9_sumout ),
	.cout(\Add11~10 ),
	.shareout(\Add11~11 ));
defparam \Add11~9 .extended_lut = "off";
defparam \Add11~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~9 .shared_arith = "on";

cyclonev_lcell_comb \Add11~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][5]~q ),
	.datad(!\butterfly_st1[2][0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~10 ),
	.sharein(\Add11~11 ),
	.combout(),
	.sumout(\Add11~13_sumout ),
	.cout(\Add11~14 ),
	.shareout(\Add11~15 ));
defparam \Add11~13 .extended_lut = "off";
defparam \Add11~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~13 .shared_arith = "on";

cyclonev_lcell_comb \Add11~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][6]~q ),
	.datad(!\butterfly_st1[2][0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~14 ),
	.sharein(\Add11~15 ),
	.combout(),
	.sumout(\Add11~17_sumout ),
	.cout(\Add11~18 ),
	.shareout(\Add11~19 ));
defparam \Add11~17 .extended_lut = "off";
defparam \Add11~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~17 .shared_arith = "on";

cyclonev_lcell_comb \Add11~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][7]~q ),
	.datad(!\butterfly_st1[2][0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~18 ),
	.sharein(\Add11~19 ),
	.combout(),
	.sumout(\Add11~21_sumout ),
	.cout(\Add11~22 ),
	.shareout(\Add11~23 ));
defparam \Add11~21 .extended_lut = "off";
defparam \Add11~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~21 .shared_arith = "on";

cyclonev_lcell_comb \Add11~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][8]~q ),
	.datad(!\butterfly_st1[2][0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~22 ),
	.sharein(\Add11~23 ),
	.combout(),
	.sumout(\Add11~25_sumout ),
	.cout(\Add11~26 ),
	.shareout(\Add11~27 ));
defparam \Add11~25 .extended_lut = "off";
defparam \Add11~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~25 .shared_arith = "on";

cyclonev_lcell_comb \Add11~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][8]~q ),
	.datad(!\butterfly_st1[2][0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~26 ),
	.sharein(\Add11~27 ),
	.combout(),
	.sumout(\Add11~29_sumout ),
	.cout(),
	.shareout());
defparam \Add11~29 .extended_lut = "off";
defparam \Add11~29 .lut_mask = 64'h0000000000000FF0;
defparam \Add11~29 .shared_arith = "on";

cyclonev_lcell_comb \Add15~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][1][2]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][0][2]~q ),
	.datag(gnd),
	.cin(\Add15~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~1_sumout ),
	.cout(\Add15~2 ),
	.shareout());
defparam \Add15~1 .extended_lut = "off";
defparam \Add15~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~1 .shared_arith = "off";

dffeas \butterfly_st2[3][1][1] (
	.clk(clk),
	.d(\Add15~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][1] .power_up = "low";

cyclonev_lcell_comb \Add15~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][1][3]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][0][3]~q ),
	.datag(gnd),
	.cin(\Add15~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~5_sumout ),
	.cout(\Add15~6 ),
	.shareout());
defparam \Add15~5 .extended_lut = "off";
defparam \Add15~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~5 .shared_arith = "off";

cyclonev_lcell_comb \Add15~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][1][4]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][0][4]~q ),
	.datag(gnd),
	.cin(\Add15~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~9_sumout ),
	.cout(\Add15~10 ),
	.shareout());
defparam \Add15~9 .extended_lut = "off";
defparam \Add15~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~9 .shared_arith = "off";

cyclonev_lcell_comb \Add15~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[3][0][5]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[2][1][5]~q ),
	.datag(gnd),
	.cin(\Add15~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~13_sumout ),
	.cout(\Add15~14 ),
	.shareout());
defparam \Add15~13 .extended_lut = "off";
defparam \Add15~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~13 .shared_arith = "off";

cyclonev_lcell_comb \Add15~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[3][0][6]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[2][1][6]~q ),
	.datag(gnd),
	.cin(\Add15~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~17_sumout ),
	.cout(\Add15~18 ),
	.shareout());
defparam \Add15~17 .extended_lut = "off";
defparam \Add15~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~17 .shared_arith = "off";

cyclonev_lcell_comb \Add15~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[3][0][7]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[2][1][7]~q ),
	.datag(gnd),
	.cin(\Add15~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~21_sumout ),
	.cout(\Add15~22 ),
	.shareout());
defparam \Add15~21 .extended_lut = "off";
defparam \Add15~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~21 .shared_arith = "off";

cyclonev_lcell_comb \Add15~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[3][0][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[2][1][8]~q ),
	.datag(gnd),
	.cin(\Add15~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~25_sumout ),
	.cout(\Add15~26 ),
	.shareout());
defparam \Add15~25 .extended_lut = "off";
defparam \Add15~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~25 .shared_arith = "off";

cyclonev_lcell_comb \Add15~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[3][0][8]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[2][1][8]~q ),
	.datag(gnd),
	.cin(\Add15~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~29_sumout ),
	.cout(),
	.shareout());
defparam \Add15~29 .extended_lut = "off";
defparam \Add15~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~29 .shared_arith = "off";

dffeas \butterfly_st1[1][0][7] (
	.clk(clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][7] .power_up = "low";

dffeas \butterfly_st1[0][0][7] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][7] .power_up = "low";

dffeas \butterfly_st1[1][1][7] (
	.clk(clk),
	.d(\Add5~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][7] .power_up = "low";

dffeas \butterfly_st1[0][1][7] (
	.clk(clk),
	.d(\Add4~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][7] .power_up = "low";

dffeas \butterfly_st1[2][0][2] (
	.clk(clk),
	.d(\Add2~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][2] .power_up = "low";

dffeas \butterfly_st1[3][1][2] (
	.clk(clk),
	.d(\Add7~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][2] .power_up = "low";

cyclonev_lcell_comb \Add9~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][1]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][1]~q ),
	.datag(gnd),
	.cin(\Add9~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~33_sumout ),
	.cout(\Add9~34 ),
	.shareout());
defparam \Add9~33 .extended_lut = "off";
defparam \Add9~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~33 .shared_arith = "off";

dffeas \butterfly_st2[1][0][0] (
	.clk(clk),
	.d(\Add9~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[1][0][0] .power_up = "low";

dffeas \butterfly_st1[2][0][3] (
	.clk(clk),
	.d(\Add2~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][3] .power_up = "low";

dffeas \butterfly_st1[3][1][3] (
	.clk(clk),
	.d(\Add7~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][3] .power_up = "low";

dffeas \butterfly_st1[2][0][4] (
	.clk(clk),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][4] .power_up = "low";

dffeas \butterfly_st1[3][1][4] (
	.clk(clk),
	.d(\Add7~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][4] .power_up = "low";

dffeas \butterfly_st1[2][0][5] (
	.clk(clk),
	.d(\Add2~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][5] .power_up = "low";

dffeas \butterfly_st1[3][1][5] (
	.clk(clk),
	.d(\Add7~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][5] .power_up = "low";

dffeas \butterfly_st1[2][0][6] (
	.clk(clk),
	.d(\Add2~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][6] .power_up = "low";

dffeas \butterfly_st1[3][1][6] (
	.clk(clk),
	.d(\Add7~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][6] .power_up = "low";

dffeas \butterfly_st1[2][0][7] (
	.clk(clk),
	.d(\Add2~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][7] .power_up = "low";

dffeas \butterfly_st1[3][1][7] (
	.clk(clk),
	.d(\Add7~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][7] .power_up = "low";

dffeas \butterfly_st1[2][0][8] (
	.clk(clk),
	.d(\Add2~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][8] .power_up = "low";

dffeas \butterfly_st1[3][1][8] (
	.clk(clk),
	.d(\Add7~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][8] .power_up = "low";

dffeas \butterfly_st1[3][0][2] (
	.clk(clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][2] .power_up = "low";

dffeas \butterfly_st1[2][1][2] (
	.clk(clk),
	.d(\Add6~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][2] .power_up = "low";

cyclonev_lcell_comb \Add13~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][0][1]~q ),
	.datad(!\butterfly_st1[2][1][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add13~38 ),
	.sharein(\Add13~39 ),
	.combout(),
	.sumout(\Add13~33_sumout ),
	.cout(\Add13~34 ),
	.shareout(\Add13~35 ));
defparam \Add13~33 .extended_lut = "off";
defparam \Add13~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add13~33 .shared_arith = "on";

dffeas \butterfly_st2[1][1][0] (
	.clk(clk),
	.d(\Add13~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[1][1][0] .power_up = "low";

dffeas \butterfly_st1[3][0][3] (
	.clk(clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][3] .power_up = "low";

dffeas \butterfly_st1[2][1][3] (
	.clk(clk),
	.d(\Add6~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][3] .power_up = "low";

dffeas \butterfly_st1[3][0][4] (
	.clk(clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][4] .power_up = "low";

dffeas \butterfly_st1[2][1][4] (
	.clk(clk),
	.d(\Add6~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][4] .power_up = "low";

dffeas \butterfly_st1[2][1][5] (
	.clk(clk),
	.d(\Add6~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][5] .power_up = "low";

dffeas \butterfly_st1[3][0][5] (
	.clk(clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][5] .power_up = "low";

dffeas \butterfly_st1[2][1][6] (
	.clk(clk),
	.d(\Add6~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][6] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][6] .power_up = "low";

dffeas \butterfly_st1[3][0][6] (
	.clk(clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][6]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][6] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][6] .power_up = "low";

dffeas \butterfly_st1[2][1][7] (
	.clk(clk),
	.d(\Add6~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][7] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][7] .power_up = "low";

dffeas \butterfly_st1[3][0][7] (
	.clk(clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][7]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][7] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][7] .power_up = "low";

dffeas \butterfly_st1[2][1][8] (
	.clk(clk),
	.d(\Add6~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][8] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][8] .power_up = "low";

dffeas \butterfly_st1[3][0][8] (
	.clk(clk),
	.d(\Add3~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][8]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][8] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][8] .power_up = "low";

dffeas \butterfly_st1[0][0][2] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][2] .power_up = "low";

dffeas \butterfly_st1[1][0][2] (
	.clk(clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][2] .power_up = "low";

cyclonev_lcell_comb \Add10~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][1]~q ),
	.datad(!\butterfly_st1[1][0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~38 ),
	.sharein(\Add10~39 ),
	.combout(),
	.sumout(\Add10~33_sumout ),
	.cout(\Add10~34 ),
	.shareout(\Add10~35 ));
defparam \Add10~33 .extended_lut = "off";
defparam \Add10~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~33 .shared_arith = "on";

dffeas \butterfly_st2[2][0][0] (
	.clk(clk),
	.d(\Add10~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[2][0][0] .power_up = "low";

dffeas \butterfly_st1[0][0][3] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][3] .power_up = "low";

dffeas \butterfly_st1[1][0][3] (
	.clk(clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][3] .power_up = "low";

dffeas \butterfly_st1[0][0][4] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][4] .power_up = "low";

dffeas \butterfly_st1[1][0][4] (
	.clk(clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][4] .power_up = "low";

dffeas \butterfly_st1[0][0][5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][5] .power_up = "low";

dffeas \butterfly_st1[1][0][5] (
	.clk(clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][5] .power_up = "low";

dffeas \butterfly_st1[0][1][2] (
	.clk(clk),
	.d(\Add4~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][2] .power_up = "low";

dffeas \butterfly_st1[1][1][2] (
	.clk(clk),
	.d(\Add5~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][2] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][2] .power_up = "low";

cyclonev_lcell_comb \Add14~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][1]~q ),
	.datad(!\butterfly_st1[1][1][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add14~38 ),
	.sharein(\Add14~39 ),
	.combout(),
	.sumout(\Add14~33_sumout ),
	.cout(\Add14~34 ),
	.shareout(\Add14~35 ));
defparam \Add14~33 .extended_lut = "off";
defparam \Add14~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~33 .shared_arith = "on";

dffeas \butterfly_st2[2][1][0] (
	.clk(clk),
	.d(\Add14~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[2][1][0] .power_up = "low";

dffeas \butterfly_st1[0][1][3] (
	.clk(clk),
	.d(\Add4~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][3] .power_up = "low";

dffeas \butterfly_st1[1][1][3] (
	.clk(clk),
	.d(\Add5~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][3] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][3] .power_up = "low";

dffeas \butterfly_st1[0][1][4] (
	.clk(clk),
	.d(\Add4~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][4] .power_up = "low";

dffeas \butterfly_st1[1][1][4] (
	.clk(clk),
	.d(\Add5~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][4]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][4] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][4] .power_up = "low";

dffeas \butterfly_st1[0][1][5] (
	.clk(clk),
	.d(\Add4~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][5] .power_up = "low";

dffeas \butterfly_st1[1][1][5] (
	.clk(clk),
	.d(\Add5~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][5]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][5] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][5] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][6]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][6]~q ),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][6]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][6]~q ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add8~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][4]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][4]~q ),
	.datag(gnd),
	.cin(\Add8~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~21_sumout ),
	.cout(\Add8~22 ),
	.shareout());
defparam \Add8~21 .extended_lut = "off";
defparam \Add8~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~21 .shared_arith = "off";

dffeas \butterfly_st2[0][0][3] (
	.clk(clk),
	.d(\Add8~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][3] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][3] .power_up = "low";

dffeas \butterfly_st2[0][0][2] (
	.clk(clk),
	.d(\Add8~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][2] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][2] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~1_sumout ),
	.cout(),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][6]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][6]~q ),
	.datag(gnd),
	.cin(\Add5~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~5_sumout ),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][6]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][6]~q ),
	.datag(gnd),
	.cin(\Add4~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add12~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][4]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][4]~q ),
	.datag(gnd),
	.cin(\Add12~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~21_sumout ),
	.cout(\Add12~22 ),
	.shareout());
defparam \Add12~21 .extended_lut = "off";
defparam \Add12~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~21 .shared_arith = "off";

dffeas \butterfly_st2[0][1][3] (
	.clk(clk),
	.d(\Add12~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][3]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][3] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][3] .power_up = "low";

dffeas \butterfly_st2[0][1][2] (
	.clk(clk),
	.d(\Add12~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][2]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][2] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][2] .power_up = "low";

cyclonev_lcell_comb \Add11~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][1]~q ),
	.datad(!\butterfly_st1[2][0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~38 ),
	.sharein(\Add11~39 ),
	.combout(),
	.sumout(\Add11~33_sumout ),
	.cout(\Add11~34 ),
	.shareout(\Add11~35 ));
defparam \Add11~33 .extended_lut = "off";
defparam \Add11~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~33 .shared_arith = "on";

dffeas \butterfly_st2[3][0][0] (
	.clk(clk),
	.d(\Add11~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[3][0][0] .power_up = "low";

cyclonev_lcell_comb \Add15~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][1][1]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][0][1]~q ),
	.datag(gnd),
	.cin(\Add15~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~33_sumout ),
	.cout(\Add15~34 ),
	.shareout());
defparam \Add15~33 .extended_lut = "off";
defparam \Add15~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~33 .shared_arith = "off";

dffeas \butterfly_st2[3][1][0] (
	.clk(clk),
	.d(\Add15~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[3][1][0] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~9_sumout ),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][2]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(\Add2~31 ),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout(\Add2~3 ));
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~1 .shared_arith = "on";

cyclonev_lcell_comb \Add7~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][2]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~30 ),
	.sharein(\Add7~31 ),
	.combout(),
	.sumout(\Add7~1_sumout ),
	.cout(\Add7~2 ),
	.shareout(\Add7~3 ));
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add7~1 .shared_arith = "on";

dffeas \butterfly_st1[2][0][1] (
	.clk(clk),
	.d(\Add2~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][1] .power_up = "low";

dffeas \butterfly_st1[3][1][1] (
	.clk(clk),
	.d(\Add7~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][1] .power_up = "low";

cyclonev_lcell_comb \Add9~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][0][0]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~37_sumout ),
	.cout(\Add9~38 ),
	.shareout());
defparam \Add9~37 .extended_lut = "off";
defparam \Add9~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~37 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[0][3]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[2][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(\Add2~3 ),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout(\Add2~7 ));
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add2~5 .shared_arith = "on";

cyclonev_lcell_comb \Add7~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[1][3]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[3][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~2 ),
	.sharein(\Add7~3 ),
	.combout(),
	.sumout(\Add7~5_sumout ),
	.cout(\Add7~6 ),
	.shareout(\Add7~7 ));
defparam \Add7~5 .extended_lut = "off";
defparam \Add7~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add7~5 .shared_arith = "on";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][4]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(\Add2~7 ),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout(\Add2~11 ));
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~9 .shared_arith = "on";

cyclonev_lcell_comb \Add7~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][4]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~6 ),
	.sharein(\Add7~7 ),
	.combout(),
	.sumout(\Add7~9_sumout ),
	.cout(\Add7~10 ),
	.shareout(\Add7~11 ));
defparam \Add7~9 .extended_lut = "off";
defparam \Add7~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add7~9 .shared_arith = "on";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][5]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(\Add2~11 ),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout(\Add2~15 ));
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~13 .shared_arith = "on";

cyclonev_lcell_comb \Add7~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][5]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~10 ),
	.sharein(\Add7~11 ),
	.combout(),
	.sumout(\Add7~13_sumout ),
	.cout(\Add7~14 ),
	.shareout(\Add7~15 ));
defparam \Add7~13 .extended_lut = "off";
defparam \Add7~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add7~13 .shared_arith = "on";

cyclonev_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][6]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(\Add2~15 ),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout(\Add2~19 ));
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~17 .shared_arith = "on";

cyclonev_lcell_comb \Add7~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][6]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~14 ),
	.sharein(\Add7~15 ),
	.combout(),
	.sumout(\Add7~17_sumout ),
	.cout(\Add7~18 ),
	.shareout(\Add7~19 ));
defparam \Add7~17 .extended_lut = "off";
defparam \Add7~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add7~17 .shared_arith = "on";

cyclonev_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(\Add2~19 ),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout(\Add2~23 ));
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~21 .shared_arith = "on";

cyclonev_lcell_comb \Add7~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~18 ),
	.sharein(\Add7~19 ),
	.combout(),
	.sumout(\Add7~21_sumout ),
	.cout(\Add7~22 ),
	.shareout(\Add7~23 ));
defparam \Add7~21 .extended_lut = "off";
defparam \Add7~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add7~21 .shared_arith = "on";

cyclonev_lcell_comb \Add2~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][7]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(\Add2~23 ),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(),
	.shareout());
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h0000000000000FF0;
defparam \Add2~25 .shared_arith = "on";

cyclonev_lcell_comb \Add7~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][7]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~22 ),
	.sharein(\Add7~23 ),
	.combout(),
	.sumout(\Add7~25_sumout ),
	.cout(),
	.shareout());
defparam \Add7~25 .extended_lut = "off";
defparam \Add7~25 .lut_mask = 64'h0000000000000FF0;
defparam \Add7~25 .shared_arith = "on";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][2]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(\Add3~31 ),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout(\Add3~3 ));
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~1 .shared_arith = "on";

cyclonev_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][2]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~30 ),
	.sharein(\Add6~31 ),
	.combout(),
	.sumout(\Add6~1_sumout ),
	.cout(\Add6~2 ),
	.shareout(\Add6~3 ));
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~1 .shared_arith = "on";

dffeas \butterfly_st1[3][0][1] (
	.clk(clk),
	.d(\Add3~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][1] .power_up = "low";

dffeas \butterfly_st1[2][1][1] (
	.clk(clk),
	.d(\Add6~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][1] .power_up = "low";

cyclonev_lcell_comb \Add13~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][0][0]~q ),
	.datad(!\butterfly_st1[2][1][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add13~37_sumout ),
	.cout(\Add13~38 ),
	.shareout(\Add13~39 ));
defparam \Add13~37 .extended_lut = "off";
defparam \Add13~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add13~37 .shared_arith = "on";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][3]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(\Add3~3 ),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout(\Add3~7 ));
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~5 .shared_arith = "on";

cyclonev_lcell_comb \Add6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[0][3]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[2][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~2 ),
	.sharein(\Add6~3 ),
	.combout(),
	.sumout(\Add6~5_sumout ),
	.cout(\Add6~6 ),
	.shareout(\Add6~7 ));
defparam \Add6~5 .extended_lut = "off";
defparam \Add6~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add6~5 .shared_arith = "on";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][4]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(\Add3~7 ),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout(\Add3~11 ));
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~9 .shared_arith = "on";

cyclonev_lcell_comb \Add6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][4]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~6 ),
	.sharein(\Add6~7 ),
	.combout(),
	.sumout(\Add6~9_sumout ),
	.cout(\Add6~10 ),
	.shareout(\Add6~11 ));
defparam \Add6~9 .extended_lut = "off";
defparam \Add6~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~9 .shared_arith = "on";

cyclonev_lcell_comb \Add6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][5]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~10 ),
	.sharein(\Add6~11 ),
	.combout(),
	.sumout(\Add6~13_sumout ),
	.cout(\Add6~14 ),
	.shareout(\Add6~15 ));
defparam \Add6~13 .extended_lut = "off";
defparam \Add6~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~13 .shared_arith = "on";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][5]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(\Add3~11 ),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout(\Add3~15 ));
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~13 .shared_arith = "on";

cyclonev_lcell_comb \Add6~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][6]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~14 ),
	.sharein(\Add6~15 ),
	.combout(),
	.sumout(\Add6~17_sumout ),
	.cout(\Add6~18 ),
	.shareout(\Add6~19 ));
defparam \Add6~17 .extended_lut = "off";
defparam \Add6~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~17 .shared_arith = "on";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][6]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(\Add3~15 ),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout(\Add3~19 ));
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~17 .shared_arith = "on";

cyclonev_lcell_comb \Add6~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~18 ),
	.sharein(\Add6~19 ),
	.combout(),
	.sumout(\Add6~21_sumout ),
	.cout(\Add6~22 ),
	.shareout(\Add6~23 ));
defparam \Add6~21 .extended_lut = "off";
defparam \Add6~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~21 .shared_arith = "on";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(\Add3~19 ),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout(\Add3~23 ));
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~21 .shared_arith = "on";

cyclonev_lcell_comb \Add6~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][7]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~22 ),
	.sharein(\Add6~23 ),
	.combout(),
	.sumout(\Add6~25_sumout ),
	.cout(),
	.shareout());
defparam \Add6~25 .extended_lut = "off";
defparam \Add6~25 .lut_mask = 64'h0000000000000FF0;
defparam \Add6~25 .shared_arith = "on";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][7]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(\Add3~23 ),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h0000000000000FF0;
defparam \Add3~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][2]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][2]~q ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][2]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][2]~q ),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~13 .shared_arith = "off";

dffeas \butterfly_st1[0][0][1] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][1] .power_up = "low";

dffeas \butterfly_st1[1][0][1] (
	.clk(clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][1] .power_up = "low";

cyclonev_lcell_comb \Add10~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][0][0]~q ),
	.datad(!\butterfly_st1[1][0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~37_sumout ),
	.cout(\Add10~38 ),
	.shareout(\Add10~39 ));
defparam \Add10~37 .extended_lut = "off";
defparam \Add10~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add10~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[2][3]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[0][3]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][3]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][3]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][4]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][4]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][4]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][4]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][5]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][5]~q ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][5]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][5]~q ),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][2]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][2]~q ),
	.datag(gnd),
	.cin(\Add4~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][2]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][2]~q ),
	.datag(gnd),
	.cin(\Add5~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~13_sumout ),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~13 .shared_arith = "off";

dffeas \butterfly_st1[0][1][1] (
	.clk(clk),
	.d(\Add4~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][1] .power_up = "low";

dffeas \butterfly_st1[1][1][1] (
	.clk(clk),
	.d(\Add5~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][1] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][1] .power_up = "low";

cyclonev_lcell_comb \Add14~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[0][1][0]~q ),
	.datad(!\butterfly_st1[1][1][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add14~37_sumout ),
	.cout(\Add14~38 ),
	.shareout(\Add14~39 ));
defparam \Add14~37 .extended_lut = "off";
defparam \Add14~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add14~37 .shared_arith = "on";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[2][3]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[0][3]~q ),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[3][3]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[1][3]~q ),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~17_sumout ),
	.cout(\Add5~18 ),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~17 .shared_arith = "off";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][4]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][4]~q ),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(\Add4~22 ),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~21 .shared_arith = "off";

cyclonev_lcell_comb \Add5~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][4]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][4]~q ),
	.datag(gnd),
	.cin(\Add5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~21_sumout ),
	.cout(\Add5~22 ),
	.shareout());
defparam \Add5~21 .extended_lut = "off";
defparam \Add5~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~21 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][5]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][5]~q ),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(\Add4~26 ),
	.shareout());
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~25 .shared_arith = "off";

cyclonev_lcell_comb \Add5~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][5]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][5]~q ),
	.datag(gnd),
	.cin(\Add5~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~25_sumout ),
	.cout(\Add5~26 ),
	.shareout());
defparam \Add5~25 .extended_lut = "off";
defparam \Add5~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~25 .shared_arith = "off";

cyclonev_lcell_comb \Add8~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][3]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][3]~q ),
	.datag(gnd),
	.cin(\Add8~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~25_sumout ),
	.cout(\Add8~26 ),
	.shareout());
defparam \Add8~25 .extended_lut = "off";
defparam \Add8~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~25 .shared_arith = "off";

cyclonev_lcell_comb \Add8~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][2]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][2]~q ),
	.datag(gnd),
	.cin(\Add8~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~29_sumout ),
	.cout(\Add8~30 ),
	.shareout());
defparam \Add8~29 .extended_lut = "off";
defparam \Add8~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~29 .shared_arith = "off";

dffeas \butterfly_st2[0][0][1] (
	.clk(clk),
	.d(\Add8~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][1] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][1] .power_up = "low";

cyclonev_lcell_comb \Add12~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][3]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][3]~q ),
	.datag(gnd),
	.cin(\Add12~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~25_sumout ),
	.cout(\Add12~26 ),
	.shareout());
defparam \Add12~25 .extended_lut = "off";
defparam \Add12~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~25 .shared_arith = "off";

cyclonev_lcell_comb \Add12~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][2]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][2]~q ),
	.datag(gnd),
	.cin(\Add12~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~29_sumout ),
	.cout(\Add12~30 ),
	.shareout());
defparam \Add12~29 .extended_lut = "off";
defparam \Add12~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~29 .shared_arith = "off";

dffeas \butterfly_st2[0][1][1] (
	.clk(clk),
	.d(\Add12~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][1]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][1] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][1] .power_up = "low";

cyclonev_lcell_comb \Add11~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\butterfly_st1[3][1][0]~q ),
	.datad(!\butterfly_st1[2][0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~37_sumout ),
	.cout(\Add11~38 ),
	.shareout(\Add11~39 ));
defparam \Add11~37 .extended_lut = "off";
defparam \Add11~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add11~37 .shared_arith = "on";

cyclonev_lcell_comb \Add15~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[2][1][0]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[3][0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~37_sumout ),
	.cout(\Add15~38 ),
	.shareout());
defparam \Add15~37 .extended_lut = "off";
defparam \Add15~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~37 .shared_arith = "off";

cyclonev_lcell_comb \Add2~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[0][1]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[2][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(\Add2~35 ),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout(\Add2~31 ));
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add2~29 .shared_arith = "on";

cyclonev_lcell_comb \Add7~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[3][1]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~34 ),
	.sharein(\Add7~35 ),
	.combout(),
	.sumout(\Add7~29_sumout ),
	.cout(\Add7~30 ),
	.shareout(\Add7~31 ));
defparam \Add7~29 .extended_lut = "off";
defparam \Add7~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add7~29 .shared_arith = "on";

dffeas \butterfly_st1[2][0][0] (
	.clk(clk),
	.d(\Add2~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][0][0] .power_up = "low";

dffeas \butterfly_st1[3][1][0] (
	.clk(clk),
	.d(\Add7~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][1][0] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][1]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(\Add3~35 ),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout(\Add3~31 ));
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~29 .shared_arith = "on";

cyclonev_lcell_comb \Add6~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][1]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~34 ),
	.sharein(\Add6~35 ),
	.combout(),
	.sumout(\Add6~29_sumout ),
	.cout(\Add6~30 ),
	.shareout(\Add6~31 ));
defparam \Add6~29 .extended_lut = "off";
defparam \Add6~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~29 .shared_arith = "on";

dffeas \butterfly_st1[3][0][0] (
	.clk(clk),
	.d(\Add3~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[3][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[3][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[3][0][0] .power_up = "low";

dffeas \butterfly_st1[2][1][0] (
	.clk(clk),
	.d(\Add6~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[2][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[2][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[2][1][0] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[2][1]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[0][1]~q ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][1]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][1]~q ),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~29 .shared_arith = "off";

dffeas \butterfly_st1[0][0][0] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][0][0] .power_up = "low";

dffeas \butterfly_st1[1][0][0] (
	.clk(clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][0][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][0][0] .power_up = "low";

cyclonev_lcell_comb \Add4~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][1]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][1]~q ),
	.datag(gnd),
	.cin(\Add4~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~29_sumout ),
	.cout(\Add4~30 ),
	.shareout());
defparam \Add4~29 .extended_lut = "off";
defparam \Add4~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~29 .shared_arith = "off";

cyclonev_lcell_comb \Add5~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[1][1]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[3][1]~q ),
	.datag(gnd),
	.cin(\Add5~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~29_sumout ),
	.cout(\Add5~30 ),
	.shareout());
defparam \Add5~29 .extended_lut = "off";
defparam \Add5~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~29 .shared_arith = "off";

dffeas \butterfly_st1[0][1][0] (
	.clk(clk),
	.d(\Add4~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[0][1][0] .power_up = "low";

dffeas \butterfly_st1[1][1][0] (
	.clk(clk),
	.d(\Add5~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st1[1][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st1[1][1][0] .is_wysiwyg = "true";
defparam \butterfly_st1[1][1][0] .power_up = "low";

cyclonev_lcell_comb \Add8~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][1]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][1]~q ),
	.datag(gnd),
	.cin(\Add8~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~33_sumout ),
	.cout(\Add8~34 ),
	.shareout());
defparam \Add8~33 .extended_lut = "off";
defparam \Add8~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~33 .shared_arith = "off";

dffeas \butterfly_st2[0][0][0] (
	.clk(clk),
	.d(\Add8~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][0][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][0][0] .is_wysiwyg = "true";
defparam \butterfly_st2[0][0][0] .power_up = "low";

cyclonev_lcell_comb \Add12~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][1]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][1]~q ),
	.datag(gnd),
	.cin(\Add12~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~33_sumout ),
	.cout(\Add12~34 ),
	.shareout());
defparam \Add12~33 .extended_lut = "off";
defparam \Add12~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~33 .shared_arith = "off";

dffeas \butterfly_st2[0][1][0] (
	.clk(clk),
	.d(\Add12~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\butterfly_st2[0][1][0]~q ),
	.prn(vcc));
defparam \butterfly_st2[0][1][0] .is_wysiwyg = "true";
defparam \butterfly_st2[0][1][0] .power_up = "low";

cyclonev_lcell_comb \Add2~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[2][0]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout(\Add2~35 ));
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add2~33 .shared_arith = "on";

cyclonev_lcell_comb \Add7~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[1][0]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[3][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~33_sumout ),
	.cout(\Add7~34 ),
	.shareout(\Add7~35 ));
defparam \Add7~33 .extended_lut = "off";
defparam \Add7~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add7~33 .shared_arith = "on";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|r_array_out[3][0]~q ),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout(\Add3~35 ));
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add3~33 .shared_arith = "on";

cyclonev_lcell_comb \Add6~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\gen_disc:bfp_scale|i_array_out[2][0]~q ),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~33_sumout ),
	.cout(\Add6~34 ),
	.shareout(\Add6~35 ));
defparam \Add6~33 .extended_lut = "off";
defparam \Add6~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add6~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[0][0]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[2][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|r_array_out[1][0]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|r_array_out[3][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~33 .shared_arith = "off";

cyclonev_lcell_comb \Add4~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[0][0]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[2][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~33_sumout ),
	.cout(\Add4~34 ),
	.shareout());
defparam \Add4~33 .extended_lut = "off";
defparam \Add4~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add4~33 .shared_arith = "off";

cyclonev_lcell_comb \Add5~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_disc:bfp_scale|i_array_out[3][0]~q ),
	.datae(gnd),
	.dataf(!\gen_disc:bfp_scale|i_array_out[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~33_sumout ),
	.cout(\Add5~34 ),
	.shareout());
defparam \Add5~33 .extended_lut = "off";
defparam \Add5~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add5~33 .shared_arith = "off";

cyclonev_lcell_comb \Add8~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][0][0]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~37_sumout ),
	.cout(\Add8~38 ),
	.shareout());
defparam \Add8~37 .extended_lut = "off";
defparam \Add8~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add8~37 .shared_arith = "off";

cyclonev_lcell_comb \Add12~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\butterfly_st1[1][1][0]~q ),
	.datae(gnd),
	.dataf(!\butterfly_st1[0][1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~37_sumout ),
	.cout(\Add12~38 ),
	.shareout());
defparam \Add12~37 .extended_lut = "off";
defparam \Add12~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add12~37 .shared_arith = "off";

dffeas \reg_no_twiddle[6][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle603),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][3] .power_up = "low";

dffeas \reg_no_twiddle[6][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle607),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][7] .power_up = "low";

dffeas \reg_no_twiddle[6][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle617),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][7] .power_up = "low";

dffeas \reg_no_twiddle[6][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle613),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][3] .power_up = "low";

dffeas \reg_no_twiddle[6][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle604),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][4] .power_up = "low";

dffeas \reg_no_twiddle[6][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle614),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][4] .power_up = "low";

dffeas \reg_no_twiddle[6][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle605),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][5] .power_up = "low";

dffeas \reg_no_twiddle[6][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle615),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][5] .power_up = "low";

dffeas \reg_no_twiddle[6][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle606),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][6] .power_up = "low";

dffeas \reg_no_twiddle[6][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle616),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][6] .power_up = "low";

dffeas \reg_no_twiddle[6][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle602),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][2] .power_up = "low";

dffeas \reg_no_twiddle[6][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle612),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][2] .power_up = "low";

dffeas \reg_no_twiddle[6][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle601),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][1] .power_up = "low";

dffeas \reg_no_twiddle[6][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle611),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][1] .power_up = "low";

dffeas \reg_no_twiddle[6][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[5][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle600),
	.prn(vcc));
defparam \reg_no_twiddle[6][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][0][0] .power_up = "low";

dffeas \reg_no_twiddle[6][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[5][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(reg_no_twiddle610),
	.prn(vcc));
defparam \reg_no_twiddle[6][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[6][1][0] .power_up = "low";

cyclonev_lcell_comb \Add16~29 (
	.dataa(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datae(gnd),
	.dataf(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~29_sumout ),
	.cout(\Add16~30 ),
	.shareout());
defparam \Add16~29 .extended_lut = "off";
defparam \Add16~29 .lut_mask = 64'h0000FF55000000FF;
defparam \Add16~29 .shared_arith = "off";

cyclonev_lcell_comb \Add16~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~25_sumout ),
	.cout(\Add16~26 ),
	.shareout());
defparam \Add16~25 .extended_lut = "off";
defparam \Add16~25 .lut_mask = 64'h00000000000000FF;
defparam \Add16~25 .shared_arith = "off";

cyclonev_lcell_comb \Add16~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~21_sumout ),
	.cout(\Add16~22 ),
	.shareout());
defparam \Add16~21 .extended_lut = "off";
defparam \Add16~21 .lut_mask = 64'h00000000000000FF;
defparam \Add16~21 .shared_arith = "off";

cyclonev_lcell_comb \Add16~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~1_sumout ),
	.cout(\Add16~2 ),
	.shareout());
defparam \Add16~1 .extended_lut = "off";
defparam \Add16~1 .lut_mask = 64'h00000000000000FF;
defparam \Add16~1 .shared_arith = "off";

dffeas \reg_no_twiddle[0][0][3] (
	.clk(clk),
	.d(\Add16~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][3] .power_up = "low";

dffeas \reg_no_twiddle[1][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][3] .power_up = "low";

dffeas \reg_no_twiddle[2][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][3] .power_up = "low";

dffeas \reg_no_twiddle[3][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][3] .power_up = "low";

dffeas \reg_no_twiddle[4][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][3] .power_up = "low";

dffeas \reg_no_twiddle[5][0][3] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][3] .power_up = "low";

cyclonev_lcell_comb \Add16~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~9_sumout ),
	.cout(\Add16~10 ),
	.shareout());
defparam \Add16~9 .extended_lut = "off";
defparam \Add16~9 .lut_mask = 64'h00000000000000FF;
defparam \Add16~9 .shared_arith = "off";

cyclonev_lcell_comb \Add16~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~13_sumout ),
	.cout(\Add16~14 ),
	.shareout());
defparam \Add16~13 .extended_lut = "off";
defparam \Add16~13 .lut_mask = 64'h00000000000000FF;
defparam \Add16~13 .shared_arith = "off";

cyclonev_lcell_comb \Add16~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~17_sumout ),
	.cout(\Add16~18 ),
	.shareout());
defparam \Add16~17 .extended_lut = "off";
defparam \Add16~17 .lut_mask = 64'h00000000000000FF;
defparam \Add16~17 .shared_arith = "off";

cyclonev_lcell_comb \Add16~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~5_sumout ),
	.cout(),
	.shareout());
defparam \Add16~5 .extended_lut = "off";
defparam \Add16~5 .lut_mask = 64'h00000000000000FF;
defparam \Add16~5 .shared_arith = "off";

dffeas \reg_no_twiddle[0][0][7] (
	.clk(clk),
	.d(\Add16~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][7] .power_up = "low";

dffeas \reg_no_twiddle[1][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][7] .power_up = "low";

dffeas \reg_no_twiddle[2][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][7] .power_up = "low";

dffeas \reg_no_twiddle[3][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][7] .power_up = "low";

dffeas \reg_no_twiddle[4][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][7] .power_up = "low";

dffeas \reg_no_twiddle[5][0][7] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][7] .power_up = "low";

cyclonev_lcell_comb \Add17~29 (
	.dataa(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datae(gnd),
	.dataf(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~29_sumout ),
	.cout(\Add17~30 ),
	.shareout());
defparam \Add17~29 .extended_lut = "off";
defparam \Add17~29 .lut_mask = 64'h0000FF55000000FF;
defparam \Add17~29 .shared_arith = "off";

cyclonev_lcell_comb \Add17~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~25_sumout ),
	.cout(\Add17~26 ),
	.shareout());
defparam \Add17~25 .extended_lut = "off";
defparam \Add17~25 .lut_mask = 64'h00000000000000FF;
defparam \Add17~25 .shared_arith = "off";

cyclonev_lcell_comb \Add17~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~21_sumout ),
	.cout(\Add17~22 ),
	.shareout());
defparam \Add17~21 .extended_lut = "off";
defparam \Add17~21 .lut_mask = 64'h00000000000000FF;
defparam \Add17~21 .shared_arith = "off";

cyclonev_lcell_comb \Add17~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~5_sumout ),
	.cout(\Add17~6 ),
	.shareout());
defparam \Add17~5 .extended_lut = "off";
defparam \Add17~5 .lut_mask = 64'h00000000000000FF;
defparam \Add17~5 .shared_arith = "off";

cyclonev_lcell_comb \Add17~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~9_sumout ),
	.cout(\Add17~10 ),
	.shareout());
defparam \Add17~9 .extended_lut = "off";
defparam \Add17~9 .lut_mask = 64'h00000000000000FF;
defparam \Add17~9 .shared_arith = "off";

cyclonev_lcell_comb \Add17~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~13_sumout ),
	.cout(\Add17~14 ),
	.shareout());
defparam \Add17~13 .extended_lut = "off";
defparam \Add17~13 .lut_mask = 64'h00000000000000FF;
defparam \Add17~13 .shared_arith = "off";

cyclonev_lcell_comb \Add17~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~17_sumout ),
	.cout(\Add17~18 ),
	.shareout());
defparam \Add17~17 .extended_lut = "off";
defparam \Add17~17 .lut_mask = 64'h00000000000000FF;
defparam \Add17~17 .shared_arith = "off";

cyclonev_lcell_comb \Add17~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~1_sumout ),
	.cout(),
	.shareout());
defparam \Add17~1 .extended_lut = "off";
defparam \Add17~1 .lut_mask = 64'h00000000000000FF;
defparam \Add17~1 .shared_arith = "off";

dffeas \reg_no_twiddle[0][1][7] (
	.clk(clk),
	.d(\Add17~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][7] .power_up = "low";

dffeas \reg_no_twiddle[1][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][7] .power_up = "low";

dffeas \reg_no_twiddle[2][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][7] .power_up = "low";

dffeas \reg_no_twiddle[3][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][7] .power_up = "low";

dffeas \reg_no_twiddle[4][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][7] .power_up = "low";

dffeas \reg_no_twiddle[5][1][7] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][7]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][7] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][7] .power_up = "low";

dffeas \reg_no_twiddle[0][1][3] (
	.clk(clk),
	.d(\Add17~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][3] .power_up = "low";

dffeas \reg_no_twiddle[1][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][3] .power_up = "low";

dffeas \reg_no_twiddle[2][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][3] .power_up = "low";

dffeas \reg_no_twiddle[3][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][3] .power_up = "low";

dffeas \reg_no_twiddle[4][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][3] .power_up = "low";

dffeas \reg_no_twiddle[5][1][3] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][3]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][3] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][3] .power_up = "low";

dffeas \reg_no_twiddle[0][0][4] (
	.clk(clk),
	.d(\Add16~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][4] .power_up = "low";

dffeas \reg_no_twiddle[1][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][4] .power_up = "low";

dffeas \reg_no_twiddle[2][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][4] .power_up = "low";

dffeas \reg_no_twiddle[3][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][4] .power_up = "low";

dffeas \reg_no_twiddle[4][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][4] .power_up = "low";

dffeas \reg_no_twiddle[5][0][4] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][4] .power_up = "low";

dffeas \reg_no_twiddle[0][1][4] (
	.clk(clk),
	.d(\Add17~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][4] .power_up = "low";

dffeas \reg_no_twiddle[1][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][4] .power_up = "low";

dffeas \reg_no_twiddle[2][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][4] .power_up = "low";

dffeas \reg_no_twiddle[3][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][4] .power_up = "low";

dffeas \reg_no_twiddle[4][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][4] .power_up = "low";

dffeas \reg_no_twiddle[5][1][4] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][4]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][4] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][4] .power_up = "low";

dffeas \reg_no_twiddle[0][0][5] (
	.clk(clk),
	.d(\Add16~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][5] .power_up = "low";

dffeas \reg_no_twiddle[1][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][5] .power_up = "low";

dffeas \reg_no_twiddle[2][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][5] .power_up = "low";

dffeas \reg_no_twiddle[3][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][5] .power_up = "low";

dffeas \reg_no_twiddle[4][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][5] .power_up = "low";

dffeas \reg_no_twiddle[5][0][5] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][5] .power_up = "low";

dffeas \reg_no_twiddle[0][1][5] (
	.clk(clk),
	.d(\Add17~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][5] .power_up = "low";

dffeas \reg_no_twiddle[1][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][5] .power_up = "low";

dffeas \reg_no_twiddle[2][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][5] .power_up = "low";

dffeas \reg_no_twiddle[3][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][5] .power_up = "low";

dffeas \reg_no_twiddle[4][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][5] .power_up = "low";

dffeas \reg_no_twiddle[5][1][5] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][5]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][5] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][5] .power_up = "low";

dffeas \reg_no_twiddle[0][0][6] (
	.clk(clk),
	.d(\Add16~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][6] .power_up = "low";

dffeas \reg_no_twiddle[1][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][6] .power_up = "low";

dffeas \reg_no_twiddle[2][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][6] .power_up = "low";

dffeas \reg_no_twiddle[3][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][6] .power_up = "low";

dffeas \reg_no_twiddle[4][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][6] .power_up = "low";

dffeas \reg_no_twiddle[5][0][6] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][6] .power_up = "low";

dffeas \reg_no_twiddle[0][1][6] (
	.clk(clk),
	.d(\Add17~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][6] .power_up = "low";

dffeas \reg_no_twiddle[1][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][6] .power_up = "low";

dffeas \reg_no_twiddle[2][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][6] .power_up = "low";

dffeas \reg_no_twiddle[3][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][6] .power_up = "low";

dffeas \reg_no_twiddle[4][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][6] .power_up = "low";

dffeas \reg_no_twiddle[5][1][6] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][6]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][6] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][6] .power_up = "low";

dffeas \reg_no_twiddle[0][0][2] (
	.clk(clk),
	.d(\Add16~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][2] .power_up = "low";

dffeas \reg_no_twiddle[1][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][2] .power_up = "low";

dffeas \reg_no_twiddle[2][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][2] .power_up = "low";

dffeas \reg_no_twiddle[3][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][2] .power_up = "low";

dffeas \reg_no_twiddle[4][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][2] .power_up = "low";

dffeas \reg_no_twiddle[5][0][2] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][2] .power_up = "low";

dffeas \reg_no_twiddle[0][1][2] (
	.clk(clk),
	.d(\Add17~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][2] .power_up = "low";

dffeas \reg_no_twiddle[1][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][2] .power_up = "low";

dffeas \reg_no_twiddle[2][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][2] .power_up = "low";

dffeas \reg_no_twiddle[3][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][2] .power_up = "low";

dffeas \reg_no_twiddle[4][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][2] .power_up = "low";

dffeas \reg_no_twiddle[5][1][2] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][2]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][2] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][2] .power_up = "low";

dffeas \reg_no_twiddle[0][0][1] (
	.clk(clk),
	.d(\Add16~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][1] .power_up = "low";

dffeas \reg_no_twiddle[1][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][1] .power_up = "low";

dffeas \reg_no_twiddle[2][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][1] .power_up = "low";

dffeas \reg_no_twiddle[3][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][1] .power_up = "low";

dffeas \reg_no_twiddle[4][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][1] .power_up = "low";

dffeas \reg_no_twiddle[5][0][1] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][1] .power_up = "low";

dffeas \reg_no_twiddle[0][1][1] (
	.clk(clk),
	.d(\Add17~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][1] .power_up = "low";

dffeas \reg_no_twiddle[1][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][1] .power_up = "low";

dffeas \reg_no_twiddle[2][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][1] .power_up = "low";

dffeas \reg_no_twiddle[3][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][1] .power_up = "low";

dffeas \reg_no_twiddle[4][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][1] .power_up = "low";

dffeas \reg_no_twiddle[5][1][1] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][1]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][1] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][1] .power_up = "low";

dffeas \reg_no_twiddle[0][0][0] (
	.clk(clk),
	.d(\Add16~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][0][0] .power_up = "low";

dffeas \reg_no_twiddle[1][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[0][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][0][0] .power_up = "low";

dffeas \reg_no_twiddle[2][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[1][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][0][0] .power_up = "low";

dffeas \reg_no_twiddle[3][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[2][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][0][0] .power_up = "low";

dffeas \reg_no_twiddle[4][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[3][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][0][0] .power_up = "low";

dffeas \reg_no_twiddle[5][0][0] (
	.clk(clk),
	.d(\reg_no_twiddle[4][0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][0][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][0][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][0][0] .power_up = "low";

dffeas \reg_no_twiddle[0][1][0] (
	.clk(clk),
	.d(\Add17~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[0][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[0][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[0][1][0] .power_up = "low";

dffeas \reg_no_twiddle[1][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[0][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[1][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[1][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[1][1][0] .power_up = "low";

dffeas \reg_no_twiddle[2][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[1][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[2][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[2][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[2][1][0] .power_up = "low";

dffeas \reg_no_twiddle[3][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[2][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[3][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[3][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[3][1][0] .power_up = "low";

dffeas \reg_no_twiddle[4][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[3][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[4][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[4][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[4][1][0] .power_up = "low";

dffeas \reg_no_twiddle[5][1][0] (
	.clk(clk),
	.d(\reg_no_twiddle[4][1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\reg_no_twiddle[5][1][0]~q ),
	.prn(vcc));
defparam \reg_no_twiddle[5][1][0] .is_wysiwyg = "true";
defparam \reg_no_twiddle[5][1][0] .power_up = "low";

endmodule

module IFFT_apn_fft_cmult_cpx2 (
	twiddle_data010,
	twiddle_data011,
	twiddle_data012,
	twiddle_data013,
	twiddle_data014,
	twiddle_data015,
	twiddle_data016,
	twiddle_data017,
	twiddle_data007,
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_3_11,
	tdl_arr_7_11,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_5_1,
	tdl_arr_5_11,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_0_1,
	tdl_arr_0_11,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	twiddle_data000,
	twiddle_data001,
	twiddle_data002,
	twiddle_data003,
	twiddle_data004,
	twiddle_data005,
	twiddle_data006,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	twiddle_data010;
input 	twiddle_data011;
input 	twiddle_data012;
input 	twiddle_data013;
input 	twiddle_data014;
input 	twiddle_data015;
input 	twiddle_data016;
input 	twiddle_data017;
input 	twiddle_data007;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_3_11;
output 	tdl_arr_7_11;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_5_1;
output 	tdl_arr_5_11;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	twiddle_data000;
input 	twiddle_data001;
input 	twiddle_data002;
input 	twiddle_data003;
input 	twiddle_data004;
input 	twiddle_data005;
input 	twiddle_data006;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \result_r_tmp[11]~q ;
wire \result_r_tmp[15]~q ;
wire \result_i_tmp[11]~q ;
wire \result_i_tmp[15]~q ;
wire \result_r_tmp[12]~q ;
wire \result_i_tmp[12]~q ;
wire \result_r_tmp[13]~q ;
wire \result_i_tmp[13]~q ;
wire \result_r_tmp[14]~q ;
wire \result_i_tmp[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ;
wire \result_r_tmp[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ;
wire \result_i_tmp[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ;
wire \result_r_tmp[9]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ;
wire \result_i_tmp[9]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ;
wire \result_r_tmp[8]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ;
wire \result_i_tmp[8]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ;
wire \result_r_tmp[7]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ;
wire \result_i_tmp[7]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ;
wire \result_r_tmp[6]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ;
wire \result_i_tmp[6]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ;
wire \result_r_tmp[5]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ;
wire \result_i_tmp[5]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ;
wire \result_r_tmp[4]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ;
wire \result_i_tmp[4]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ;
wire \result_r_tmp[3]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ;
wire \result_i_tmp[3]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ;
wire \result_r_tmp[2]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ;
wire \result_i_tmp[2]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ;
wire \result_r_tmp[1]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ;
wire \result_i_tmp[1]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ;
wire \result_r_tmp[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ;
wire \result_i_tmp[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ;


IFFT_asj_fft_pround u0(
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_11(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_r_tmp_11(\result_r_tmp[11]~q ),
	.result_r_tmp_15(\result_r_tmp[15]~q ),
	.result_r_tmp_12(\result_r_tmp[12]~q ),
	.result_r_tmp_13(\result_r_tmp[13]~q ),
	.result_r_tmp_14(\result_r_tmp[14]~q ),
	.result_r_tmp_10(\result_r_tmp[10]~q ),
	.result_r_tmp_9(\result_r_tmp[9]~q ),
	.pipeline_dffe_10(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.result_r_tmp_8(\result_r_tmp[8]~q ),
	.pipeline_dffe_9(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.result_r_tmp_7(\result_r_tmp[7]~q ),
	.pipeline_dffe_8(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.result_r_tmp_6(\result_r_tmp[6]~q ),
	.result_r_tmp_5(\result_r_tmp[5]~q ),
	.result_r_tmp_4(\result_r_tmp[4]~q ),
	.result_r_tmp_3(\result_r_tmp[3]~q ),
	.result_r_tmp_2(\result_r_tmp[2]~q ),
	.result_r_tmp_1(\result_r_tmp[1]~q ),
	.result_r_tmp_0(\result_r_tmp[0]~q ),
	.clk(clk));

IFFT_apn_fft_mult_cpx \gen_infr_4cpx:calc_mult_4cpx (
	.d({twiddle_data017,twiddle_data016,twiddle_data015,twiddle_data014,twiddle_data013,twiddle_data012,twiddle_data011,twiddle_data010}),
	.c({twiddle_data007,twiddle_data006,twiddle_data005,twiddle_data004,twiddle_data003,twiddle_data002,twiddle_data001,twiddle_data000}),
	.global_clock_enable(global_clock_enable),
	.rout_sig2_11(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ),
	.rout_sig2_15(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ),
	.iout_sig2_11(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ),
	.iout_sig2_15(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ),
	.rout_sig2_12(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ),
	.iout_sig2_12(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ),
	.rout_sig2_13(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ),
	.iout_sig2_13(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ),
	.rout_sig2_14(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ),
	.iout_sig2_14(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ),
	.rout_sig2_10(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ),
	.iout_sig2_10(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ),
	.rout_sig2_9(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ),
	.iout_sig2_9(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ),
	.rout_sig2_8(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ),
	.iout_sig2_8(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ),
	.b({pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.a({pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.rout_sig2_7(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ),
	.iout_sig2_7(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ),
	.rout_sig2_6(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ),
	.iout_sig2_6(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ),
	.rout_sig2_5(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ),
	.iout_sig2_5(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ),
	.rout_sig2_4(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ),
	.iout_sig2_4(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ),
	.rout_sig2_3(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ),
	.iout_sig2_3(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ),
	.rout_sig2_2(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ),
	.iout_sig2_2(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ),
	.rout_sig2_1(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ),
	.iout_sig2_1(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ),
	.rout_sig2_0(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ),
	.iout_sig2_0(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ),
	.clk(clk),
	.reset(reset));

IFFT_asj_fft_tdl imag_delay(
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_6_1(tdl_arr_6_11),
	.data_in({\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,
\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ,
\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q }),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_0_1(tdl_arr_0_1),
	.clk(clk));

IFFT_asj_fft_tdl_1 real_delay(
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_6_1(tdl_arr_6_1),
	.data_in({\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,
\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ,
\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q }),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_0_1(tdl_arr_0_11),
	.clk(clk));

IFFT_asj_fft_pround_1 u1(
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_11(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_i_tmp_11(\result_i_tmp[11]~q ),
	.result_i_tmp_15(\result_i_tmp[15]~q ),
	.result_i_tmp_12(\result_i_tmp[12]~q ),
	.result_i_tmp_13(\result_i_tmp[13]~q ),
	.result_i_tmp_14(\result_i_tmp[14]~q ),
	.result_i_tmp_10(\result_i_tmp[10]~q ),
	.result_i_tmp_9(\result_i_tmp[9]~q ),
	.pipeline_dffe_10(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.result_i_tmp_8(\result_i_tmp[8]~q ),
	.pipeline_dffe_9(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.result_i_tmp_7(\result_i_tmp[7]~q ),
	.pipeline_dffe_8(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.result_i_tmp_6(\result_i_tmp[6]~q ),
	.result_i_tmp_5(\result_i_tmp[5]~q ),
	.result_i_tmp_4(\result_i_tmp[4]~q ),
	.result_i_tmp_3(\result_i_tmp[3]~q ),
	.result_i_tmp_2(\result_i_tmp[2]~q ),
	.result_i_tmp_1(\result_i_tmp[1]~q ),
	.result_i_tmp_0(\result_i_tmp[0]~q ),
	.clk(clk));

dffeas \result_r_tmp[11] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[11]~q ),
	.prn(vcc));
defparam \result_r_tmp[11] .is_wysiwyg = "true";
defparam \result_r_tmp[11] .power_up = "low";

dffeas \result_r_tmp[15] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[15]~q ),
	.prn(vcc));
defparam \result_r_tmp[15] .is_wysiwyg = "true";
defparam \result_r_tmp[15] .power_up = "low";

dffeas \result_i_tmp[11] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[11]~q ),
	.prn(vcc));
defparam \result_i_tmp[11] .is_wysiwyg = "true";
defparam \result_i_tmp[11] .power_up = "low";

dffeas \result_i_tmp[15] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[15]~q ),
	.prn(vcc));
defparam \result_i_tmp[15] .is_wysiwyg = "true";
defparam \result_i_tmp[15] .power_up = "low";

dffeas \result_r_tmp[12] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[12]~q ),
	.prn(vcc));
defparam \result_r_tmp[12] .is_wysiwyg = "true";
defparam \result_r_tmp[12] .power_up = "low";

dffeas \result_i_tmp[12] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[12]~q ),
	.prn(vcc));
defparam \result_i_tmp[12] .is_wysiwyg = "true";
defparam \result_i_tmp[12] .power_up = "low";

dffeas \result_r_tmp[13] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[13]~q ),
	.prn(vcc));
defparam \result_r_tmp[13] .is_wysiwyg = "true";
defparam \result_r_tmp[13] .power_up = "low";

dffeas \result_i_tmp[13] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[13]~q ),
	.prn(vcc));
defparam \result_i_tmp[13] .is_wysiwyg = "true";
defparam \result_i_tmp[13] .power_up = "low";

dffeas \result_r_tmp[14] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[14]~q ),
	.prn(vcc));
defparam \result_r_tmp[14] .is_wysiwyg = "true";
defparam \result_r_tmp[14] .power_up = "low";

dffeas \result_i_tmp[14] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[14]~q ),
	.prn(vcc));
defparam \result_i_tmp[14] .is_wysiwyg = "true";
defparam \result_i_tmp[14] .power_up = "low";

dffeas \result_r_tmp[10] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[10]~q ),
	.prn(vcc));
defparam \result_r_tmp[10] .is_wysiwyg = "true";
defparam \result_r_tmp[10] .power_up = "low";

dffeas \result_i_tmp[10] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[10]~q ),
	.prn(vcc));
defparam \result_i_tmp[10] .is_wysiwyg = "true";
defparam \result_i_tmp[10] .power_up = "low";

dffeas \result_r_tmp[9] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[9]~q ),
	.prn(vcc));
defparam \result_r_tmp[9] .is_wysiwyg = "true";
defparam \result_r_tmp[9] .power_up = "low";

dffeas \result_i_tmp[9] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[9]~q ),
	.prn(vcc));
defparam \result_i_tmp[9] .is_wysiwyg = "true";
defparam \result_i_tmp[9] .power_up = "low";

dffeas \result_r_tmp[8] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[8]~q ),
	.prn(vcc));
defparam \result_r_tmp[8] .is_wysiwyg = "true";
defparam \result_r_tmp[8] .power_up = "low";

dffeas \result_i_tmp[8] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[8]~q ),
	.prn(vcc));
defparam \result_i_tmp[8] .is_wysiwyg = "true";
defparam \result_i_tmp[8] .power_up = "low";

dffeas \result_r_tmp[7] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[7]~q ),
	.prn(vcc));
defparam \result_r_tmp[7] .is_wysiwyg = "true";
defparam \result_r_tmp[7] .power_up = "low";

dffeas \result_i_tmp[7] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[7]~q ),
	.prn(vcc));
defparam \result_i_tmp[7] .is_wysiwyg = "true";
defparam \result_i_tmp[7] .power_up = "low";

dffeas \result_r_tmp[6] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[6]~q ),
	.prn(vcc));
defparam \result_r_tmp[6] .is_wysiwyg = "true";
defparam \result_r_tmp[6] .power_up = "low";

dffeas \result_i_tmp[6] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[6]~q ),
	.prn(vcc));
defparam \result_i_tmp[6] .is_wysiwyg = "true";
defparam \result_i_tmp[6] .power_up = "low";

dffeas \result_r_tmp[5] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[5]~q ),
	.prn(vcc));
defparam \result_r_tmp[5] .is_wysiwyg = "true";
defparam \result_r_tmp[5] .power_up = "low";

dffeas \result_i_tmp[5] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[5]~q ),
	.prn(vcc));
defparam \result_i_tmp[5] .is_wysiwyg = "true";
defparam \result_i_tmp[5] .power_up = "low";

dffeas \result_r_tmp[4] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[4]~q ),
	.prn(vcc));
defparam \result_r_tmp[4] .is_wysiwyg = "true";
defparam \result_r_tmp[4] .power_up = "low";

dffeas \result_i_tmp[4] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[4]~q ),
	.prn(vcc));
defparam \result_i_tmp[4] .is_wysiwyg = "true";
defparam \result_i_tmp[4] .power_up = "low";

dffeas \result_r_tmp[3] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[3]~q ),
	.prn(vcc));
defparam \result_r_tmp[3] .is_wysiwyg = "true";
defparam \result_r_tmp[3] .power_up = "low";

dffeas \result_i_tmp[3] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[3]~q ),
	.prn(vcc));
defparam \result_i_tmp[3] .is_wysiwyg = "true";
defparam \result_i_tmp[3] .power_up = "low";

dffeas \result_r_tmp[2] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[2]~q ),
	.prn(vcc));
defparam \result_r_tmp[2] .is_wysiwyg = "true";
defparam \result_r_tmp[2] .power_up = "low";

dffeas \result_i_tmp[2] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[2]~q ),
	.prn(vcc));
defparam \result_i_tmp[2] .is_wysiwyg = "true";
defparam \result_i_tmp[2] .power_up = "low";

dffeas \result_r_tmp[1] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[1]~q ),
	.prn(vcc));
defparam \result_r_tmp[1] .is_wysiwyg = "true";
defparam \result_r_tmp[1] .power_up = "low";

dffeas \result_i_tmp[1] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[1]~q ),
	.prn(vcc));
defparam \result_i_tmp[1] .is_wysiwyg = "true";
defparam \result_i_tmp[1] .power_up = "low";

dffeas \result_r_tmp[0] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[0]~q ),
	.prn(vcc));
defparam \result_r_tmp[0] .is_wysiwyg = "true";
defparam \result_r_tmp[0] .power_up = "low";

dffeas \result_i_tmp[0] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[0]~q ),
	.prn(vcc));
defparam \result_i_tmp[0] .is_wysiwyg = "true";
defparam \result_i_tmp[0] .power_up = "low";

endmodule

module IFFT_apn_fft_mult_cpx (
	d,
	c,
	global_clock_enable,
	rout_sig2_11,
	rout_sig2_15,
	iout_sig2_11,
	iout_sig2_15,
	rout_sig2_12,
	iout_sig2_12,
	rout_sig2_13,
	iout_sig2_13,
	rout_sig2_14,
	iout_sig2_14,
	rout_sig2_10,
	iout_sig2_10,
	rout_sig2_9,
	iout_sig2_9,
	rout_sig2_8,
	iout_sig2_8,
	b,
	a,
	rout_sig2_7,
	iout_sig2_7,
	rout_sig2_6,
	iout_sig2_6,
	rout_sig2_5,
	iout_sig2_5,
	rout_sig2_4,
	iout_sig2_4,
	rout_sig2_3,
	iout_sig2_3,
	rout_sig2_2,
	iout_sig2_2,
	rout_sig2_1,
	iout_sig2_1,
	rout_sig2_0,
	iout_sig2_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[7:0] d;
input 	[7:0] c;
input 	global_clock_enable;
output 	rout_sig2_11;
output 	rout_sig2_15;
output 	iout_sig2_11;
output 	iout_sig2_15;
output 	rout_sig2_12;
output 	iout_sig2_12;
output 	rout_sig2_13;
output 	iout_sig2_13;
output 	rout_sig2_14;
output 	iout_sig2_14;
output 	rout_sig2_10;
output 	iout_sig2_10;
output 	rout_sig2_9;
output 	iout_sig2_9;
output 	rout_sig2_8;
output 	iout_sig2_8;
input 	[7:0] b;
input 	[7:0] a;
output 	rout_sig2_7;
output 	iout_sig2_7;
output 	rout_sig2_6;
output 	iout_sig2_6;
output 	rout_sig2_5;
output 	iout_sig2_5;
output 	rout_sig2_4;
output 	iout_sig2_4;
output 	rout_sig2_3;
output 	iout_sig2_3;
output 	rout_sig2_2;
output 	iout_sig2_2;
output 	rout_sig2_1;
output 	iout_sig2_1;
output 	rout_sig2_0;
output 	iout_sig2_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~24 ;
wire \Add0~25 ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~28 ;
wire \Add0~29 ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~32 ;
wire \Add0~33 ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~36 ;
wire \Add0~37 ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~40 ;
wire \Add0~41 ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~44 ;
wire \Add0~45 ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~48 ;
wire \Add0~49 ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~52 ;
wire \Add0~53 ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~56 ;
wire \Add0~57 ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~60 ;
wire \Add0~61 ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~64 ;
wire \Add0~65 ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~68 ;
wire \Add0~69 ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \Add1~24 ;
wire \Add1~25 ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~28 ;
wire \Add1~29 ;
wire \Add1~30 ;
wire \Add1~31 ;
wire \Add1~32 ;
wire \Add1~33 ;
wire \Add1~34 ;
wire \Add1~35 ;
wire \Add1~36 ;
wire \Add1~37 ;
wire \Add1~38 ;
wire \Add1~39 ;
wire \Add1~40 ;
wire \Add1~41 ;
wire \Add1~42 ;
wire \Add1~43 ;
wire \Add1~44 ;
wire \Add1~45 ;
wire \Add1~46 ;
wire \Add1~47 ;
wire \Add1~48 ;
wire \Add1~49 ;
wire \Add1~50 ;
wire \Add1~51 ;
wire \Add1~52 ;
wire \Add1~53 ;
wire \Add1~54 ;
wire \Add1~55 ;
wire \Add1~56 ;
wire \Add1~57 ;
wire \Add1~58 ;
wire \Add1~59 ;
wire \Add1~60 ;
wire \Add1~61 ;
wire \Add1~62 ;
wire \Add1~63 ;
wire \Add1~64 ;
wire \Add1~65 ;
wire \Add1~66 ;
wire \Add1~67 ;
wire \Add1~68 ;
wire \Add1~69 ;
wire \Add1~70 ;
wire \Add1~71 ;
wire \d_reg[0]~q ;
wire \d_reg[1]~q ;
wire \d_reg[2]~q ;
wire \d_reg[3]~q ;
wire \d_reg[4]~q ;
wire \d_reg[5]~q ;
wire \d_reg[6]~q ;
wire \d_reg[7]~q ;
wire \b_reg[0]~q ;
wire \b_reg[1]~q ;
wire \b_reg[2]~q ;
wire \b_reg[3]~q ;
wire \b_reg[4]~q ;
wire \b_reg[5]~q ;
wire \b_reg[6]~q ;
wire \b_reg[7]~q ;
wire \c_reg[0]~q ;
wire \c_reg[1]~q ;
wire \c_reg[2]~q ;
wire \c_reg[3]~q ;
wire \c_reg[4]~q ;
wire \c_reg[5]~q ;
wire \c_reg[6]~q ;
wire \c_reg[7]~q ;
wire \a_reg[0]~q ;
wire \a_reg[1]~q ;
wire \a_reg[2]~q ;
wire \a_reg[3]~q ;
wire \a_reg[4]~q ;
wire \a_reg[5]~q ;
wire \a_reg[6]~q ;
wire \a_reg[7]~q ;
wire \Add0~19 ;
wire \rout_sig[11]~q ;
wire \Add0~23 ;
wire \rout_sig[15]~q ;
wire \Add1~19 ;
wire \iout_sig[11]~q ;
wire \Add1~23 ;
wire \iout_sig[15]~q ;
wire \Add0~20 ;
wire \rout_sig[12]~q ;
wire \Add1~20 ;
wire \iout_sig[12]~q ;
wire \Add0~21 ;
wire \rout_sig[13]~q ;
wire \Add1~21 ;
wire \iout_sig[13]~q ;
wire \Add0~22 ;
wire \rout_sig[14]~q ;
wire \Add1~22 ;
wire \iout_sig[14]~q ;
wire \Add0~18 ;
wire \rout_sig[10]~q ;
wire \Add1~18 ;
wire \iout_sig[10]~q ;
wire \Add0~17 ;
wire \rout_sig[9]~q ;
wire \Add1~17 ;
wire \iout_sig[9]~q ;
wire \Add0~16 ;
wire \rout_sig[8]~q ;
wire \Add1~16 ;
wire \iout_sig[8]~q ;
wire \Add0~15 ;
wire \rout_sig[7]~q ;
wire \Add1~15 ;
wire \iout_sig[7]~q ;
wire \Add0~14 ;
wire \rout_sig[6]~q ;
wire \Add1~14 ;
wire \iout_sig[6]~q ;
wire \Add0~13 ;
wire \rout_sig[5]~q ;
wire \Add1~13 ;
wire \iout_sig[5]~q ;
wire \Add0~12 ;
wire \rout_sig[4]~q ;
wire \Add1~12 ;
wire \iout_sig[4]~q ;
wire \Add0~11 ;
wire \rout_sig[3]~q ;
wire \Add1~11 ;
wire \iout_sig[3]~q ;
wire \Add0~10 ;
wire \rout_sig[2]~q ;
wire \Add1~10 ;
wire \iout_sig[2]~q ;
wire \Add0~9 ;
wire \rout_sig[1]~q ;
wire \Add1~9 ;
wire \iout_sig[1]~q ;
wire \Add0~8_resulta ;
wire \rout_sig[0]~q ;
wire \Add1~8_resulta ;
wire \iout_sig[0]~q ;

wire [63:0] \Add0~8_RESULTA_bus ;
wire [63:0] \Add1~8_RESULTA_bus ;

assign \Add0~8_resulta  = \Add0~8_RESULTA_bus [0];
assign \Add0~9  = \Add0~8_RESULTA_bus [1];
assign \Add0~10  = \Add0~8_RESULTA_bus [2];
assign \Add0~11  = \Add0~8_RESULTA_bus [3];
assign \Add0~12  = \Add0~8_RESULTA_bus [4];
assign \Add0~13  = \Add0~8_RESULTA_bus [5];
assign \Add0~14  = \Add0~8_RESULTA_bus [6];
assign \Add0~15  = \Add0~8_RESULTA_bus [7];
assign \Add0~16  = \Add0~8_RESULTA_bus [8];
assign \Add0~17  = \Add0~8_RESULTA_bus [9];
assign \Add0~18  = \Add0~8_RESULTA_bus [10];
assign \Add0~19  = \Add0~8_RESULTA_bus [11];
assign \Add0~20  = \Add0~8_RESULTA_bus [12];
assign \Add0~21  = \Add0~8_RESULTA_bus [13];
assign \Add0~22  = \Add0~8_RESULTA_bus [14];
assign \Add0~23  = \Add0~8_RESULTA_bus [15];
assign \Add0~24  = \Add0~8_RESULTA_bus [16];
assign \Add0~25  = \Add0~8_RESULTA_bus [17];
assign \Add0~26  = \Add0~8_RESULTA_bus [18];
assign \Add0~27  = \Add0~8_RESULTA_bus [19];
assign \Add0~28  = \Add0~8_RESULTA_bus [20];
assign \Add0~29  = \Add0~8_RESULTA_bus [21];
assign \Add0~30  = \Add0~8_RESULTA_bus [22];
assign \Add0~31  = \Add0~8_RESULTA_bus [23];
assign \Add0~32  = \Add0~8_RESULTA_bus [24];
assign \Add0~33  = \Add0~8_RESULTA_bus [25];
assign \Add0~34  = \Add0~8_RESULTA_bus [26];
assign \Add0~35  = \Add0~8_RESULTA_bus [27];
assign \Add0~36  = \Add0~8_RESULTA_bus [28];
assign \Add0~37  = \Add0~8_RESULTA_bus [29];
assign \Add0~38  = \Add0~8_RESULTA_bus [30];
assign \Add0~39  = \Add0~8_RESULTA_bus [31];
assign \Add0~40  = \Add0~8_RESULTA_bus [32];
assign \Add0~41  = \Add0~8_RESULTA_bus [33];
assign \Add0~42  = \Add0~8_RESULTA_bus [34];
assign \Add0~43  = \Add0~8_RESULTA_bus [35];
assign \Add0~44  = \Add0~8_RESULTA_bus [36];
assign \Add0~45  = \Add0~8_RESULTA_bus [37];
assign \Add0~46  = \Add0~8_RESULTA_bus [38];
assign \Add0~47  = \Add0~8_RESULTA_bus [39];
assign \Add0~48  = \Add0~8_RESULTA_bus [40];
assign \Add0~49  = \Add0~8_RESULTA_bus [41];
assign \Add0~50  = \Add0~8_RESULTA_bus [42];
assign \Add0~51  = \Add0~8_RESULTA_bus [43];
assign \Add0~52  = \Add0~8_RESULTA_bus [44];
assign \Add0~53  = \Add0~8_RESULTA_bus [45];
assign \Add0~54  = \Add0~8_RESULTA_bus [46];
assign \Add0~55  = \Add0~8_RESULTA_bus [47];
assign \Add0~56  = \Add0~8_RESULTA_bus [48];
assign \Add0~57  = \Add0~8_RESULTA_bus [49];
assign \Add0~58  = \Add0~8_RESULTA_bus [50];
assign \Add0~59  = \Add0~8_RESULTA_bus [51];
assign \Add0~60  = \Add0~8_RESULTA_bus [52];
assign \Add0~61  = \Add0~8_RESULTA_bus [53];
assign \Add0~62  = \Add0~8_RESULTA_bus [54];
assign \Add0~63  = \Add0~8_RESULTA_bus [55];
assign \Add0~64  = \Add0~8_RESULTA_bus [56];
assign \Add0~65  = \Add0~8_RESULTA_bus [57];
assign \Add0~66  = \Add0~8_RESULTA_bus [58];
assign \Add0~67  = \Add0~8_RESULTA_bus [59];
assign \Add0~68  = \Add0~8_RESULTA_bus [60];
assign \Add0~69  = \Add0~8_RESULTA_bus [61];
assign \Add0~70  = \Add0~8_RESULTA_bus [62];
assign \Add0~71  = \Add0~8_RESULTA_bus [63];

assign \Add1~8_resulta  = \Add1~8_RESULTA_bus [0];
assign \Add1~9  = \Add1~8_RESULTA_bus [1];
assign \Add1~10  = \Add1~8_RESULTA_bus [2];
assign \Add1~11  = \Add1~8_RESULTA_bus [3];
assign \Add1~12  = \Add1~8_RESULTA_bus [4];
assign \Add1~13  = \Add1~8_RESULTA_bus [5];
assign \Add1~14  = \Add1~8_RESULTA_bus [6];
assign \Add1~15  = \Add1~8_RESULTA_bus [7];
assign \Add1~16  = \Add1~8_RESULTA_bus [8];
assign \Add1~17  = \Add1~8_RESULTA_bus [9];
assign \Add1~18  = \Add1~8_RESULTA_bus [10];
assign \Add1~19  = \Add1~8_RESULTA_bus [11];
assign \Add1~20  = \Add1~8_RESULTA_bus [12];
assign \Add1~21  = \Add1~8_RESULTA_bus [13];
assign \Add1~22  = \Add1~8_RESULTA_bus [14];
assign \Add1~23  = \Add1~8_RESULTA_bus [15];
assign \Add1~24  = \Add1~8_RESULTA_bus [16];
assign \Add1~25  = \Add1~8_RESULTA_bus [17];
assign \Add1~26  = \Add1~8_RESULTA_bus [18];
assign \Add1~27  = \Add1~8_RESULTA_bus [19];
assign \Add1~28  = \Add1~8_RESULTA_bus [20];
assign \Add1~29  = \Add1~8_RESULTA_bus [21];
assign \Add1~30  = \Add1~8_RESULTA_bus [22];
assign \Add1~31  = \Add1~8_RESULTA_bus [23];
assign \Add1~32  = \Add1~8_RESULTA_bus [24];
assign \Add1~33  = \Add1~8_RESULTA_bus [25];
assign \Add1~34  = \Add1~8_RESULTA_bus [26];
assign \Add1~35  = \Add1~8_RESULTA_bus [27];
assign \Add1~36  = \Add1~8_RESULTA_bus [28];
assign \Add1~37  = \Add1~8_RESULTA_bus [29];
assign \Add1~38  = \Add1~8_RESULTA_bus [30];
assign \Add1~39  = \Add1~8_RESULTA_bus [31];
assign \Add1~40  = \Add1~8_RESULTA_bus [32];
assign \Add1~41  = \Add1~8_RESULTA_bus [33];
assign \Add1~42  = \Add1~8_RESULTA_bus [34];
assign \Add1~43  = \Add1~8_RESULTA_bus [35];
assign \Add1~44  = \Add1~8_RESULTA_bus [36];
assign \Add1~45  = \Add1~8_RESULTA_bus [37];
assign \Add1~46  = \Add1~8_RESULTA_bus [38];
assign \Add1~47  = \Add1~8_RESULTA_bus [39];
assign \Add1~48  = \Add1~8_RESULTA_bus [40];
assign \Add1~49  = \Add1~8_RESULTA_bus [41];
assign \Add1~50  = \Add1~8_RESULTA_bus [42];
assign \Add1~51  = \Add1~8_RESULTA_bus [43];
assign \Add1~52  = \Add1~8_RESULTA_bus [44];
assign \Add1~53  = \Add1~8_RESULTA_bus [45];
assign \Add1~54  = \Add1~8_RESULTA_bus [46];
assign \Add1~55  = \Add1~8_RESULTA_bus [47];
assign \Add1~56  = \Add1~8_RESULTA_bus [48];
assign \Add1~57  = \Add1~8_RESULTA_bus [49];
assign \Add1~58  = \Add1~8_RESULTA_bus [50];
assign \Add1~59  = \Add1~8_RESULTA_bus [51];
assign \Add1~60  = \Add1~8_RESULTA_bus [52];
assign \Add1~61  = \Add1~8_RESULTA_bus [53];
assign \Add1~62  = \Add1~8_RESULTA_bus [54];
assign \Add1~63  = \Add1~8_RESULTA_bus [55];
assign \Add1~64  = \Add1~8_RESULTA_bus [56];
assign \Add1~65  = \Add1~8_RESULTA_bus [57];
assign \Add1~66  = \Add1~8_RESULTA_bus [58];
assign \Add1~67  = \Add1~8_RESULTA_bus [59];
assign \Add1~68  = \Add1~8_RESULTA_bus [60];
assign \Add1~69  = \Add1~8_RESULTA_bus [61];
assign \Add1~70  = \Add1~8_RESULTA_bus [62];
assign \Add1~71  = \Add1~8_RESULTA_bus [63];

dffeas \rout_sig2[11] (
	.clk(clk),
	.d(\rout_sig[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_11),
	.prn(vcc));
defparam \rout_sig2[11] .is_wysiwyg = "true";
defparam \rout_sig2[11] .power_up = "low";

dffeas \rout_sig2[15] (
	.clk(clk),
	.d(\rout_sig[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_15),
	.prn(vcc));
defparam \rout_sig2[15] .is_wysiwyg = "true";
defparam \rout_sig2[15] .power_up = "low";

dffeas \iout_sig2[11] (
	.clk(clk),
	.d(\iout_sig[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_11),
	.prn(vcc));
defparam \iout_sig2[11] .is_wysiwyg = "true";
defparam \iout_sig2[11] .power_up = "low";

dffeas \iout_sig2[15] (
	.clk(clk),
	.d(\iout_sig[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_15),
	.prn(vcc));
defparam \iout_sig2[15] .is_wysiwyg = "true";
defparam \iout_sig2[15] .power_up = "low";

dffeas \rout_sig2[12] (
	.clk(clk),
	.d(\rout_sig[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_12),
	.prn(vcc));
defparam \rout_sig2[12] .is_wysiwyg = "true";
defparam \rout_sig2[12] .power_up = "low";

dffeas \iout_sig2[12] (
	.clk(clk),
	.d(\iout_sig[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_12),
	.prn(vcc));
defparam \iout_sig2[12] .is_wysiwyg = "true";
defparam \iout_sig2[12] .power_up = "low";

dffeas \rout_sig2[13] (
	.clk(clk),
	.d(\rout_sig[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_13),
	.prn(vcc));
defparam \rout_sig2[13] .is_wysiwyg = "true";
defparam \rout_sig2[13] .power_up = "low";

dffeas \iout_sig2[13] (
	.clk(clk),
	.d(\iout_sig[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_13),
	.prn(vcc));
defparam \iout_sig2[13] .is_wysiwyg = "true";
defparam \iout_sig2[13] .power_up = "low";

dffeas \rout_sig2[14] (
	.clk(clk),
	.d(\rout_sig[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_14),
	.prn(vcc));
defparam \rout_sig2[14] .is_wysiwyg = "true";
defparam \rout_sig2[14] .power_up = "low";

dffeas \iout_sig2[14] (
	.clk(clk),
	.d(\iout_sig[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_14),
	.prn(vcc));
defparam \iout_sig2[14] .is_wysiwyg = "true";
defparam \iout_sig2[14] .power_up = "low";

dffeas \rout_sig2[10] (
	.clk(clk),
	.d(\rout_sig[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_10),
	.prn(vcc));
defparam \rout_sig2[10] .is_wysiwyg = "true";
defparam \rout_sig2[10] .power_up = "low";

dffeas \iout_sig2[10] (
	.clk(clk),
	.d(\iout_sig[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_10),
	.prn(vcc));
defparam \iout_sig2[10] .is_wysiwyg = "true";
defparam \iout_sig2[10] .power_up = "low";

dffeas \rout_sig2[9] (
	.clk(clk),
	.d(\rout_sig[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_9),
	.prn(vcc));
defparam \rout_sig2[9] .is_wysiwyg = "true";
defparam \rout_sig2[9] .power_up = "low";

dffeas \iout_sig2[9] (
	.clk(clk),
	.d(\iout_sig[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_9),
	.prn(vcc));
defparam \iout_sig2[9] .is_wysiwyg = "true";
defparam \iout_sig2[9] .power_up = "low";

dffeas \rout_sig2[8] (
	.clk(clk),
	.d(\rout_sig[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_8),
	.prn(vcc));
defparam \rout_sig2[8] .is_wysiwyg = "true";
defparam \rout_sig2[8] .power_up = "low";

dffeas \iout_sig2[8] (
	.clk(clk),
	.d(\iout_sig[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_8),
	.prn(vcc));
defparam \iout_sig2[8] .is_wysiwyg = "true";
defparam \iout_sig2[8] .power_up = "low";

dffeas \rout_sig2[7] (
	.clk(clk),
	.d(\rout_sig[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_7),
	.prn(vcc));
defparam \rout_sig2[7] .is_wysiwyg = "true";
defparam \rout_sig2[7] .power_up = "low";

dffeas \iout_sig2[7] (
	.clk(clk),
	.d(\iout_sig[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_7),
	.prn(vcc));
defparam \iout_sig2[7] .is_wysiwyg = "true";
defparam \iout_sig2[7] .power_up = "low";

dffeas \rout_sig2[6] (
	.clk(clk),
	.d(\rout_sig[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_6),
	.prn(vcc));
defparam \rout_sig2[6] .is_wysiwyg = "true";
defparam \rout_sig2[6] .power_up = "low";

dffeas \iout_sig2[6] (
	.clk(clk),
	.d(\iout_sig[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_6),
	.prn(vcc));
defparam \iout_sig2[6] .is_wysiwyg = "true";
defparam \iout_sig2[6] .power_up = "low";

dffeas \rout_sig2[5] (
	.clk(clk),
	.d(\rout_sig[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_5),
	.prn(vcc));
defparam \rout_sig2[5] .is_wysiwyg = "true";
defparam \rout_sig2[5] .power_up = "low";

dffeas \iout_sig2[5] (
	.clk(clk),
	.d(\iout_sig[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_5),
	.prn(vcc));
defparam \iout_sig2[5] .is_wysiwyg = "true";
defparam \iout_sig2[5] .power_up = "low";

dffeas \rout_sig2[4] (
	.clk(clk),
	.d(\rout_sig[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_4),
	.prn(vcc));
defparam \rout_sig2[4] .is_wysiwyg = "true";
defparam \rout_sig2[4] .power_up = "low";

dffeas \iout_sig2[4] (
	.clk(clk),
	.d(\iout_sig[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_4),
	.prn(vcc));
defparam \iout_sig2[4] .is_wysiwyg = "true";
defparam \iout_sig2[4] .power_up = "low";

dffeas \rout_sig2[3] (
	.clk(clk),
	.d(\rout_sig[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_3),
	.prn(vcc));
defparam \rout_sig2[3] .is_wysiwyg = "true";
defparam \rout_sig2[3] .power_up = "low";

dffeas \iout_sig2[3] (
	.clk(clk),
	.d(\iout_sig[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_3),
	.prn(vcc));
defparam \iout_sig2[3] .is_wysiwyg = "true";
defparam \iout_sig2[3] .power_up = "low";

dffeas \rout_sig2[2] (
	.clk(clk),
	.d(\rout_sig[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_2),
	.prn(vcc));
defparam \rout_sig2[2] .is_wysiwyg = "true";
defparam \rout_sig2[2] .power_up = "low";

dffeas \iout_sig2[2] (
	.clk(clk),
	.d(\iout_sig[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_2),
	.prn(vcc));
defparam \iout_sig2[2] .is_wysiwyg = "true";
defparam \iout_sig2[2] .power_up = "low";

dffeas \rout_sig2[1] (
	.clk(clk),
	.d(\rout_sig[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_1),
	.prn(vcc));
defparam \rout_sig2[1] .is_wysiwyg = "true";
defparam \rout_sig2[1] .power_up = "low";

dffeas \iout_sig2[1] (
	.clk(clk),
	.d(\iout_sig[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_1),
	.prn(vcc));
defparam \iout_sig2[1] .is_wysiwyg = "true";
defparam \iout_sig2[1] .power_up = "low";

dffeas \rout_sig2[0] (
	.clk(clk),
	.d(\rout_sig[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_0),
	.prn(vcc));
defparam \rout_sig2[0] .is_wysiwyg = "true";
defparam \rout_sig2[0] .power_up = "low";

dffeas \iout_sig2[0] (
	.clk(clk),
	.d(\iout_sig[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_0),
	.prn(vcc));
defparam \iout_sig2[0] .is_wysiwyg = "true";
defparam \iout_sig2[0] .power_up = "low";

dffeas \d_reg[0] (
	.clk(clk),
	.d(d[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[0]~q ),
	.prn(vcc));
defparam \d_reg[0] .is_wysiwyg = "true";
defparam \d_reg[0] .power_up = "low";

dffeas \d_reg[1] (
	.clk(clk),
	.d(d[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[1]~q ),
	.prn(vcc));
defparam \d_reg[1] .is_wysiwyg = "true";
defparam \d_reg[1] .power_up = "low";

dffeas \d_reg[2] (
	.clk(clk),
	.d(d[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[2]~q ),
	.prn(vcc));
defparam \d_reg[2] .is_wysiwyg = "true";
defparam \d_reg[2] .power_up = "low";

dffeas \d_reg[3] (
	.clk(clk),
	.d(d[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[3]~q ),
	.prn(vcc));
defparam \d_reg[3] .is_wysiwyg = "true";
defparam \d_reg[3] .power_up = "low";

dffeas \d_reg[4] (
	.clk(clk),
	.d(d[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[4]~q ),
	.prn(vcc));
defparam \d_reg[4] .is_wysiwyg = "true";
defparam \d_reg[4] .power_up = "low";

dffeas \d_reg[5] (
	.clk(clk),
	.d(d[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[5]~q ),
	.prn(vcc));
defparam \d_reg[5] .is_wysiwyg = "true";
defparam \d_reg[5] .power_up = "low";

dffeas \d_reg[6] (
	.clk(clk),
	.d(d[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[6]~q ),
	.prn(vcc));
defparam \d_reg[6] .is_wysiwyg = "true";
defparam \d_reg[6] .power_up = "low";

dffeas \d_reg[7] (
	.clk(clk),
	.d(d[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[7]~q ),
	.prn(vcc));
defparam \d_reg[7] .is_wysiwyg = "true";
defparam \d_reg[7] .power_up = "low";

dffeas \b_reg[0] (
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[0]~q ),
	.prn(vcc));
defparam \b_reg[0] .is_wysiwyg = "true";
defparam \b_reg[0] .power_up = "low";

dffeas \b_reg[1] (
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[1]~q ),
	.prn(vcc));
defparam \b_reg[1] .is_wysiwyg = "true";
defparam \b_reg[1] .power_up = "low";

dffeas \b_reg[2] (
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[2]~q ),
	.prn(vcc));
defparam \b_reg[2] .is_wysiwyg = "true";
defparam \b_reg[2] .power_up = "low";

dffeas \b_reg[3] (
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[3]~q ),
	.prn(vcc));
defparam \b_reg[3] .is_wysiwyg = "true";
defparam \b_reg[3] .power_up = "low";

dffeas \b_reg[4] (
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[4]~q ),
	.prn(vcc));
defparam \b_reg[4] .is_wysiwyg = "true";
defparam \b_reg[4] .power_up = "low";

dffeas \b_reg[5] (
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[5]~q ),
	.prn(vcc));
defparam \b_reg[5] .is_wysiwyg = "true";
defparam \b_reg[5] .power_up = "low";

dffeas \b_reg[6] (
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[6]~q ),
	.prn(vcc));
defparam \b_reg[6] .is_wysiwyg = "true";
defparam \b_reg[6] .power_up = "low";

dffeas \b_reg[7] (
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[7]~q ),
	.prn(vcc));
defparam \b_reg[7] .is_wysiwyg = "true";
defparam \b_reg[7] .power_up = "low";

dffeas \c_reg[0] (
	.clk(clk),
	.d(c[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[0]~q ),
	.prn(vcc));
defparam \c_reg[0] .is_wysiwyg = "true";
defparam \c_reg[0] .power_up = "low";

dffeas \c_reg[1] (
	.clk(clk),
	.d(c[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[1]~q ),
	.prn(vcc));
defparam \c_reg[1] .is_wysiwyg = "true";
defparam \c_reg[1] .power_up = "low";

dffeas \c_reg[2] (
	.clk(clk),
	.d(c[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[2]~q ),
	.prn(vcc));
defparam \c_reg[2] .is_wysiwyg = "true";
defparam \c_reg[2] .power_up = "low";

dffeas \c_reg[3] (
	.clk(clk),
	.d(c[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[3]~q ),
	.prn(vcc));
defparam \c_reg[3] .is_wysiwyg = "true";
defparam \c_reg[3] .power_up = "low";

dffeas \c_reg[4] (
	.clk(clk),
	.d(c[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[4]~q ),
	.prn(vcc));
defparam \c_reg[4] .is_wysiwyg = "true";
defparam \c_reg[4] .power_up = "low";

dffeas \c_reg[5] (
	.clk(clk),
	.d(c[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[5]~q ),
	.prn(vcc));
defparam \c_reg[5] .is_wysiwyg = "true";
defparam \c_reg[5] .power_up = "low";

dffeas \c_reg[6] (
	.clk(clk),
	.d(c[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[6]~q ),
	.prn(vcc));
defparam \c_reg[6] .is_wysiwyg = "true";
defparam \c_reg[6] .power_up = "low";

dffeas \c_reg[7] (
	.clk(clk),
	.d(c[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[7]~q ),
	.prn(vcc));
defparam \c_reg[7] .is_wysiwyg = "true";
defparam \c_reg[7] .power_up = "low";

dffeas \a_reg[0] (
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[0]~q ),
	.prn(vcc));
defparam \a_reg[0] .is_wysiwyg = "true";
defparam \a_reg[0] .power_up = "low";

dffeas \a_reg[1] (
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[1]~q ),
	.prn(vcc));
defparam \a_reg[1] .is_wysiwyg = "true";
defparam \a_reg[1] .power_up = "low";

dffeas \a_reg[2] (
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[2]~q ),
	.prn(vcc));
defparam \a_reg[2] .is_wysiwyg = "true";
defparam \a_reg[2] .power_up = "low";

dffeas \a_reg[3] (
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[3]~q ),
	.prn(vcc));
defparam \a_reg[3] .is_wysiwyg = "true";
defparam \a_reg[3] .power_up = "low";

dffeas \a_reg[4] (
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[4]~q ),
	.prn(vcc));
defparam \a_reg[4] .is_wysiwyg = "true";
defparam \a_reg[4] .power_up = "low";

dffeas \a_reg[5] (
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[5]~q ),
	.prn(vcc));
defparam \a_reg[5] .is_wysiwyg = "true";
defparam \a_reg[5] .power_up = "low";

dffeas \a_reg[6] (
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[6]~q ),
	.prn(vcc));
defparam \a_reg[6] .is_wysiwyg = "true";
defparam \a_reg[6] .power_up = "low";

dffeas \a_reg[7] (
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[7]~q ),
	.prn(vcc));
defparam \a_reg[7] .is_wysiwyg = "true";
defparam \a_reg[7] .power_up = "low";

cyclonev_mac \Add0~8 (
	.sub(vcc),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_reg[7]~q ,\d_reg[6]~q ,\d_reg[5]~q ,\d_reg[4]~q ,\d_reg[3]~q ,\d_reg[2]~q ,\d_reg[1]~q ,\d_reg[0]~q }),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\b_reg[7]~q ,\b_reg[6]~q ,\b_reg[5]~q ,\b_reg[4]~q ,\b_reg[3]~q ,\b_reg[2]~q ,\b_reg[1]~q ,\b_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\c_reg[7]~q ,\c_reg[6]~q ,\c_reg[5]~q ,\c_reg[4]~q ,\c_reg[3]~q ,\c_reg[2]~q ,\c_reg[1]~q ,\c_reg[0]~q }),
	.by({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\a_reg[7]~q ,\a_reg[6]~q ,\a_reg[5]~q ,\a_reg[4]~q ,\a_reg[3]~q ,\a_reg[2]~q ,\a_reg[1]~q ,\a_reg[0]~q }),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Add0~8_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Add0~8 .accumulate_clock = "none";
defparam \Add0~8 .ax_clock = "none";
defparam \Add0~8 .ax_width = 8;
defparam \Add0~8 .ay_scan_in_clock = "none";
defparam \Add0~8 .ay_scan_in_width = 8;
defparam \Add0~8 .ay_use_scan_in = "false";
defparam \Add0~8 .az_clock = "none";
defparam \Add0~8 .bx_clock = "none";
defparam \Add0~8 .bx_width = 8;
defparam \Add0~8 .by_clock = "none";
defparam \Add0~8 .by_use_scan_in = "false";
defparam \Add0~8 .by_width = 8;
defparam \Add0~8 .bz_clock = "none";
defparam \Add0~8 .coef_a_0 = 0;
defparam \Add0~8 .coef_a_1 = 0;
defparam \Add0~8 .coef_a_2 = 0;
defparam \Add0~8 .coef_a_3 = 0;
defparam \Add0~8 .coef_a_4 = 0;
defparam \Add0~8 .coef_a_5 = 0;
defparam \Add0~8 .coef_a_6 = 0;
defparam \Add0~8 .coef_a_7 = 0;
defparam \Add0~8 .coef_b_0 = 0;
defparam \Add0~8 .coef_b_1 = 0;
defparam \Add0~8 .coef_b_2 = 0;
defparam \Add0~8 .coef_b_3 = 0;
defparam \Add0~8 .coef_b_4 = 0;
defparam \Add0~8 .coef_b_5 = 0;
defparam \Add0~8 .coef_b_6 = 0;
defparam \Add0~8 .coef_b_7 = 0;
defparam \Add0~8 .coef_sel_a_clock = "none";
defparam \Add0~8 .coef_sel_b_clock = "none";
defparam \Add0~8 .delay_scan_out_ay = "false";
defparam \Add0~8 .delay_scan_out_by = "false";
defparam \Add0~8 .enable_double_accum = "false";
defparam \Add0~8 .load_const_clock = "none";
defparam \Add0~8 .load_const_value = 0;
defparam \Add0~8 .mode_sub_location = 0;
defparam \Add0~8 .negate_clock = "none";
defparam \Add0~8 .operand_source_max = "input";
defparam \Add0~8 .operand_source_may = "input";
defparam \Add0~8 .operand_source_mbx = "input";
defparam \Add0~8 .operand_source_mby = "input";
defparam \Add0~8 .operation_mode = "m18x18_sumof2";
defparam \Add0~8 .output_clock = "none";
defparam \Add0~8 .preadder_subtract_a = "false";
defparam \Add0~8 .preadder_subtract_b = "false";
defparam \Add0~8 .result_a_width = 64;
defparam \Add0~8 .signed_max = "true";
defparam \Add0~8 .signed_may = "true";
defparam \Add0~8 .signed_mbx = "true";
defparam \Add0~8 .signed_mby = "true";
defparam \Add0~8 .sub_clock = "none";
defparam \Add0~8 .use_chainadder = "false";

dffeas \rout_sig[11] (
	.clk(clk),
	.d(\Add0~19 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[11]~q ),
	.prn(vcc));
defparam \rout_sig[11] .is_wysiwyg = "true";
defparam \rout_sig[11] .power_up = "low";

dffeas \rout_sig[15] (
	.clk(clk),
	.d(\Add0~23 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[15]~q ),
	.prn(vcc));
defparam \rout_sig[15] .is_wysiwyg = "true";
defparam \rout_sig[15] .power_up = "low";

cyclonev_mac \Add1~8 (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\c_reg[7]~q ,\c_reg[6]~q ,\c_reg[5]~q ,\c_reg[4]~q ,\c_reg[3]~q ,\c_reg[2]~q ,\c_reg[1]~q ,\c_reg[0]~q }),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\b_reg[7]~q ,\b_reg[6]~q ,\b_reg[5]~q ,\b_reg[4]~q ,\b_reg[3]~q ,\b_reg[2]~q ,\b_reg[1]~q ,\b_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_reg[7]~q ,\d_reg[6]~q ,\d_reg[5]~q ,\d_reg[4]~q ,\d_reg[3]~q ,\d_reg[2]~q ,\d_reg[1]~q ,\d_reg[0]~q }),
	.by({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\a_reg[7]~q ,\a_reg[6]~q ,\a_reg[5]~q ,\a_reg[4]~q ,\a_reg[3]~q ,\a_reg[2]~q ,\a_reg[1]~q ,\a_reg[0]~q }),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Add1~8_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Add1~8 .accumulate_clock = "none";
defparam \Add1~8 .ax_clock = "none";
defparam \Add1~8 .ax_width = 8;
defparam \Add1~8 .ay_scan_in_clock = "none";
defparam \Add1~8 .ay_scan_in_width = 8;
defparam \Add1~8 .ay_use_scan_in = "false";
defparam \Add1~8 .az_clock = "none";
defparam \Add1~8 .bx_clock = "none";
defparam \Add1~8 .bx_width = 8;
defparam \Add1~8 .by_clock = "none";
defparam \Add1~8 .by_use_scan_in = "false";
defparam \Add1~8 .by_width = 8;
defparam \Add1~8 .bz_clock = "none";
defparam \Add1~8 .coef_a_0 = 0;
defparam \Add1~8 .coef_a_1 = 0;
defparam \Add1~8 .coef_a_2 = 0;
defparam \Add1~8 .coef_a_3 = 0;
defparam \Add1~8 .coef_a_4 = 0;
defparam \Add1~8 .coef_a_5 = 0;
defparam \Add1~8 .coef_a_6 = 0;
defparam \Add1~8 .coef_a_7 = 0;
defparam \Add1~8 .coef_b_0 = 0;
defparam \Add1~8 .coef_b_1 = 0;
defparam \Add1~8 .coef_b_2 = 0;
defparam \Add1~8 .coef_b_3 = 0;
defparam \Add1~8 .coef_b_4 = 0;
defparam \Add1~8 .coef_b_5 = 0;
defparam \Add1~8 .coef_b_6 = 0;
defparam \Add1~8 .coef_b_7 = 0;
defparam \Add1~8 .coef_sel_a_clock = "none";
defparam \Add1~8 .coef_sel_b_clock = "none";
defparam \Add1~8 .delay_scan_out_ay = "false";
defparam \Add1~8 .delay_scan_out_by = "false";
defparam \Add1~8 .enable_double_accum = "false";
defparam \Add1~8 .load_const_clock = "none";
defparam \Add1~8 .load_const_value = 0;
defparam \Add1~8 .mode_sub_location = 0;
defparam \Add1~8 .negate_clock = "none";
defparam \Add1~8 .operand_source_max = "input";
defparam \Add1~8 .operand_source_may = "input";
defparam \Add1~8 .operand_source_mbx = "input";
defparam \Add1~8 .operand_source_mby = "input";
defparam \Add1~8 .operation_mode = "m18x18_sumof2";
defparam \Add1~8 .output_clock = "none";
defparam \Add1~8 .preadder_subtract_a = "false";
defparam \Add1~8 .preadder_subtract_b = "false";
defparam \Add1~8 .result_a_width = 64;
defparam \Add1~8 .signed_max = "true";
defparam \Add1~8 .signed_may = "true";
defparam \Add1~8 .signed_mbx = "true";
defparam \Add1~8 .signed_mby = "true";
defparam \Add1~8 .sub_clock = "none";
defparam \Add1~8 .use_chainadder = "false";

dffeas \iout_sig[11] (
	.clk(clk),
	.d(\Add1~19 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[11]~q ),
	.prn(vcc));
defparam \iout_sig[11] .is_wysiwyg = "true";
defparam \iout_sig[11] .power_up = "low";

dffeas \iout_sig[15] (
	.clk(clk),
	.d(\Add1~23 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[15]~q ),
	.prn(vcc));
defparam \iout_sig[15] .is_wysiwyg = "true";
defparam \iout_sig[15] .power_up = "low";

dffeas \rout_sig[12] (
	.clk(clk),
	.d(\Add0~20 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[12]~q ),
	.prn(vcc));
defparam \rout_sig[12] .is_wysiwyg = "true";
defparam \rout_sig[12] .power_up = "low";

dffeas \iout_sig[12] (
	.clk(clk),
	.d(\Add1~20 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[12]~q ),
	.prn(vcc));
defparam \iout_sig[12] .is_wysiwyg = "true";
defparam \iout_sig[12] .power_up = "low";

dffeas \rout_sig[13] (
	.clk(clk),
	.d(\Add0~21 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[13]~q ),
	.prn(vcc));
defparam \rout_sig[13] .is_wysiwyg = "true";
defparam \rout_sig[13] .power_up = "low";

dffeas \iout_sig[13] (
	.clk(clk),
	.d(\Add1~21 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[13]~q ),
	.prn(vcc));
defparam \iout_sig[13] .is_wysiwyg = "true";
defparam \iout_sig[13] .power_up = "low";

dffeas \rout_sig[14] (
	.clk(clk),
	.d(\Add0~22 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[14]~q ),
	.prn(vcc));
defparam \rout_sig[14] .is_wysiwyg = "true";
defparam \rout_sig[14] .power_up = "low";

dffeas \iout_sig[14] (
	.clk(clk),
	.d(\Add1~22 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[14]~q ),
	.prn(vcc));
defparam \iout_sig[14] .is_wysiwyg = "true";
defparam \iout_sig[14] .power_up = "low";

dffeas \rout_sig[10] (
	.clk(clk),
	.d(\Add0~18 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[10]~q ),
	.prn(vcc));
defparam \rout_sig[10] .is_wysiwyg = "true";
defparam \rout_sig[10] .power_up = "low";

dffeas \iout_sig[10] (
	.clk(clk),
	.d(\Add1~18 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[10]~q ),
	.prn(vcc));
defparam \iout_sig[10] .is_wysiwyg = "true";
defparam \iout_sig[10] .power_up = "low";

dffeas \rout_sig[9] (
	.clk(clk),
	.d(\Add0~17 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[9]~q ),
	.prn(vcc));
defparam \rout_sig[9] .is_wysiwyg = "true";
defparam \rout_sig[9] .power_up = "low";

dffeas \iout_sig[9] (
	.clk(clk),
	.d(\Add1~17 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[9]~q ),
	.prn(vcc));
defparam \iout_sig[9] .is_wysiwyg = "true";
defparam \iout_sig[9] .power_up = "low";

dffeas \rout_sig[8] (
	.clk(clk),
	.d(\Add0~16 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[8]~q ),
	.prn(vcc));
defparam \rout_sig[8] .is_wysiwyg = "true";
defparam \rout_sig[8] .power_up = "low";

dffeas \iout_sig[8] (
	.clk(clk),
	.d(\Add1~16 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[8]~q ),
	.prn(vcc));
defparam \iout_sig[8] .is_wysiwyg = "true";
defparam \iout_sig[8] .power_up = "low";

dffeas \rout_sig[7] (
	.clk(clk),
	.d(\Add0~15 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[7]~q ),
	.prn(vcc));
defparam \rout_sig[7] .is_wysiwyg = "true";
defparam \rout_sig[7] .power_up = "low";

dffeas \iout_sig[7] (
	.clk(clk),
	.d(\Add1~15 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[7]~q ),
	.prn(vcc));
defparam \iout_sig[7] .is_wysiwyg = "true";
defparam \iout_sig[7] .power_up = "low";

dffeas \rout_sig[6] (
	.clk(clk),
	.d(\Add0~14 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[6]~q ),
	.prn(vcc));
defparam \rout_sig[6] .is_wysiwyg = "true";
defparam \rout_sig[6] .power_up = "low";

dffeas \iout_sig[6] (
	.clk(clk),
	.d(\Add1~14 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[6]~q ),
	.prn(vcc));
defparam \iout_sig[6] .is_wysiwyg = "true";
defparam \iout_sig[6] .power_up = "low";

dffeas \rout_sig[5] (
	.clk(clk),
	.d(\Add0~13 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[5]~q ),
	.prn(vcc));
defparam \rout_sig[5] .is_wysiwyg = "true";
defparam \rout_sig[5] .power_up = "low";

dffeas \iout_sig[5] (
	.clk(clk),
	.d(\Add1~13 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[5]~q ),
	.prn(vcc));
defparam \iout_sig[5] .is_wysiwyg = "true";
defparam \iout_sig[5] .power_up = "low";

dffeas \rout_sig[4] (
	.clk(clk),
	.d(\Add0~12 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[4]~q ),
	.prn(vcc));
defparam \rout_sig[4] .is_wysiwyg = "true";
defparam \rout_sig[4] .power_up = "low";

dffeas \iout_sig[4] (
	.clk(clk),
	.d(\Add1~12 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[4]~q ),
	.prn(vcc));
defparam \iout_sig[4] .is_wysiwyg = "true";
defparam \iout_sig[4] .power_up = "low";

dffeas \rout_sig[3] (
	.clk(clk),
	.d(\Add0~11 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[3]~q ),
	.prn(vcc));
defparam \rout_sig[3] .is_wysiwyg = "true";
defparam \rout_sig[3] .power_up = "low";

dffeas \iout_sig[3] (
	.clk(clk),
	.d(\Add1~11 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[3]~q ),
	.prn(vcc));
defparam \iout_sig[3] .is_wysiwyg = "true";
defparam \iout_sig[3] .power_up = "low";

dffeas \rout_sig[2] (
	.clk(clk),
	.d(\Add0~10 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[2]~q ),
	.prn(vcc));
defparam \rout_sig[2] .is_wysiwyg = "true";
defparam \rout_sig[2] .power_up = "low";

dffeas \iout_sig[2] (
	.clk(clk),
	.d(\Add1~10 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[2]~q ),
	.prn(vcc));
defparam \iout_sig[2] .is_wysiwyg = "true";
defparam \iout_sig[2] .power_up = "low";

dffeas \rout_sig[1] (
	.clk(clk),
	.d(\Add0~9 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[1]~q ),
	.prn(vcc));
defparam \rout_sig[1] .is_wysiwyg = "true";
defparam \rout_sig[1] .power_up = "low";

dffeas \iout_sig[1] (
	.clk(clk),
	.d(\Add1~9 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[1]~q ),
	.prn(vcc));
defparam \iout_sig[1] .is_wysiwyg = "true";
defparam \iout_sig[1] .power_up = "low";

dffeas \rout_sig[0] (
	.clk(clk),
	.d(\Add0~8_resulta ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[0]~q ),
	.prn(vcc));
defparam \rout_sig[0] .is_wysiwyg = "true";
defparam \rout_sig[0] .power_up = "low";

dffeas \iout_sig[0] (
	.clk(clk),
	.d(\Add1~8_resulta ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[0]~q ),
	.prn(vcc));
defparam \iout_sig[0] .is_wysiwyg = "true";
defparam \iout_sig[0] .power_up = "low";

endmodule

module IFFT_asj_fft_pround (
	global_clock_enable,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_1 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_r_tmp_8(result_r_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_r_tmp_7(result_r_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_1 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_8gj auto_generated(
	.clken(clken),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_r_tmp_8(result_r_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_r_tmp_7(result_r_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.clock(clock));

endmodule

module IFFT_add_sub_8gj (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_1 (
	global_clock_enable,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_2 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_i_tmp_8(result_i_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_i_tmp_7(result_i_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_2 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_8gj_1 auto_generated(
	.clken(clken),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_i_tmp_8(result_i_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_i_tmp_7(result_i_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.clock(clock));

endmodule

module IFFT_add_sub_8gj_1 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm1|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl (
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_4_1,
	tdl_arr_5_1,
	tdl_arr_6_1,
	data_in,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_4_1;
output 	tdl_arr_5_1;
output 	tdl_arr_6_1;
input 	[7:0] data_in;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][3]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;


dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_1 (
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_4_1,
	tdl_arr_5_1,
	tdl_arr_6_1,
	data_in,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_4_1;
output 	tdl_arr_5_1;
output 	tdl_arr_6_1;
input 	[7:0] data_in;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][3]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;


dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

endmodule

module IFFT_apn_fft_cmult_cpx2_1 (
	twiddle_data107,
	twiddle_data110,
	twiddle_data111,
	twiddle_data112,
	twiddle_data113,
	twiddle_data114,
	twiddle_data115,
	twiddle_data116,
	twiddle_data117,
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_3_11,
	tdl_arr_7_11,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_5_1,
	tdl_arr_5_11,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_0_1,
	tdl_arr_0_11,
	twiddle_data100,
	twiddle_data101,
	twiddle_data102,
	twiddle_data103,
	twiddle_data104,
	twiddle_data105,
	twiddle_data106,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	twiddle_data107;
input 	twiddle_data110;
input 	twiddle_data111;
input 	twiddle_data112;
input 	twiddle_data113;
input 	twiddle_data114;
input 	twiddle_data115;
input 	twiddle_data116;
input 	twiddle_data117;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_3_11;
output 	tdl_arr_7_11;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_5_1;
output 	tdl_arr_5_11;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
input 	twiddle_data100;
input 	twiddle_data101;
input 	twiddle_data102;
input 	twiddle_data103;
input 	twiddle_data104;
input 	twiddle_data105;
input 	twiddle_data106;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \result_i_tmp[11]~q ;
wire \result_i_tmp[15]~q ;
wire \result_r_tmp[11]~q ;
wire \result_r_tmp[15]~q ;
wire \result_i_tmp[12]~q ;
wire \result_r_tmp[12]~q ;
wire \result_i_tmp[13]~q ;
wire \result_r_tmp[13]~q ;
wire \result_i_tmp[14]~q ;
wire \result_r_tmp[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ;
wire \result_i_tmp[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ;
wire \result_r_tmp[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ;
wire \result_i_tmp[9]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ;
wire \result_r_tmp[9]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ;
wire \result_i_tmp[8]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ;
wire \result_r_tmp[8]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ;
wire \result_i_tmp[7]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ;
wire \result_r_tmp[7]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ;
wire \result_i_tmp[6]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ;
wire \result_r_tmp[6]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ;
wire \result_i_tmp[5]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ;
wire \result_r_tmp[5]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ;
wire \result_i_tmp[4]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ;
wire \result_r_tmp[4]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ;
wire \result_i_tmp[3]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ;
wire \result_r_tmp[3]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ;
wire \result_i_tmp[2]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ;
wire \result_r_tmp[2]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ;
wire \result_i_tmp[1]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ;
wire \result_r_tmp[1]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ;
wire \result_i_tmp[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ;
wire \result_r_tmp[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ;


IFFT_asj_fft_tdl_2 imag_delay(
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_6_1(tdl_arr_6_1),
	.data_in({\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,
\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ,
\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q }),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_0_1(tdl_arr_0_1),
	.clk(clk));

IFFT_asj_fft_tdl_3 real_delay(
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_6_1(tdl_arr_6_11),
	.data_in({\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,
\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ,
\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q }),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_0_1(tdl_arr_0_11),
	.clk(clk));

IFFT_asj_fft_pround_3 u1(
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_11(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_i_tmp_11(\result_i_tmp[11]~q ),
	.result_i_tmp_15(\result_i_tmp[15]~q ),
	.result_i_tmp_12(\result_i_tmp[12]~q ),
	.result_i_tmp_13(\result_i_tmp[13]~q ),
	.result_i_tmp_14(\result_i_tmp[14]~q ),
	.result_i_tmp_10(\result_i_tmp[10]~q ),
	.result_i_tmp_9(\result_i_tmp[9]~q ),
	.pipeline_dffe_10(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.result_i_tmp_8(\result_i_tmp[8]~q ),
	.pipeline_dffe_9(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.result_i_tmp_7(\result_i_tmp[7]~q ),
	.pipeline_dffe_8(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.result_i_tmp_6(\result_i_tmp[6]~q ),
	.result_i_tmp_5(\result_i_tmp[5]~q ),
	.result_i_tmp_4(\result_i_tmp[4]~q ),
	.result_i_tmp_3(\result_i_tmp[3]~q ),
	.result_i_tmp_2(\result_i_tmp[2]~q ),
	.result_i_tmp_1(\result_i_tmp[1]~q ),
	.result_i_tmp_0(\result_i_tmp[0]~q ),
	.clk(clk));

IFFT_asj_fft_pround_2 u0(
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_11(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_r_tmp_11(\result_r_tmp[11]~q ),
	.result_r_tmp_15(\result_r_tmp[15]~q ),
	.result_r_tmp_12(\result_r_tmp[12]~q ),
	.result_r_tmp_13(\result_r_tmp[13]~q ),
	.result_r_tmp_14(\result_r_tmp[14]~q ),
	.result_r_tmp_10(\result_r_tmp[10]~q ),
	.result_r_tmp_9(\result_r_tmp[9]~q ),
	.pipeline_dffe_10(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.result_r_tmp_8(\result_r_tmp[8]~q ),
	.pipeline_dffe_9(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.result_r_tmp_7(\result_r_tmp[7]~q ),
	.pipeline_dffe_8(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.result_r_tmp_6(\result_r_tmp[6]~q ),
	.result_r_tmp_5(\result_r_tmp[5]~q ),
	.result_r_tmp_4(\result_r_tmp[4]~q ),
	.result_r_tmp_3(\result_r_tmp[3]~q ),
	.result_r_tmp_2(\result_r_tmp[2]~q ),
	.result_r_tmp_1(\result_r_tmp[1]~q ),
	.result_r_tmp_0(\result_r_tmp[0]~q ),
	.clk(clk));

IFFT_apn_fft_mult_cpx_1 \gen_infr_4cpx:calc_mult_4cpx (
	.c({twiddle_data107,twiddle_data106,twiddle_data105,twiddle_data104,twiddle_data103,twiddle_data102,twiddle_data101,twiddle_data100}),
	.d({twiddle_data117,twiddle_data116,twiddle_data115,twiddle_data114,twiddle_data113,twiddle_data112,twiddle_data111,twiddle_data110}),
	.global_clock_enable(global_clock_enable),
	.iout_sig2_11(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ),
	.iout_sig2_15(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ),
	.rout_sig2_11(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ),
	.rout_sig2_15(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ),
	.iout_sig2_12(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ),
	.rout_sig2_12(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ),
	.iout_sig2_13(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ),
	.rout_sig2_13(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ),
	.iout_sig2_14(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ),
	.rout_sig2_14(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ),
	.iout_sig2_10(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ),
	.rout_sig2_10(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ),
	.iout_sig2_9(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ),
	.rout_sig2_9(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ),
	.iout_sig2_8(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ),
	.rout_sig2_8(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ),
	.b({pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.a({pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.iout_sig2_7(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ),
	.rout_sig2_7(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ),
	.iout_sig2_6(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ),
	.rout_sig2_6(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ),
	.iout_sig2_5(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ),
	.rout_sig2_5(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ),
	.iout_sig2_4(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ),
	.rout_sig2_4(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ),
	.iout_sig2_3(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ),
	.rout_sig2_3(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ),
	.iout_sig2_2(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ),
	.rout_sig2_2(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ),
	.iout_sig2_1(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ),
	.rout_sig2_1(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ),
	.iout_sig2_0(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ),
	.rout_sig2_0(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ),
	.clk(clk),
	.reset(reset));

dffeas \result_i_tmp[11] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[11]~q ),
	.prn(vcc));
defparam \result_i_tmp[11] .is_wysiwyg = "true";
defparam \result_i_tmp[11] .power_up = "low";

dffeas \result_i_tmp[15] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[15]~q ),
	.prn(vcc));
defparam \result_i_tmp[15] .is_wysiwyg = "true";
defparam \result_i_tmp[15] .power_up = "low";

dffeas \result_r_tmp[11] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[11]~q ),
	.prn(vcc));
defparam \result_r_tmp[11] .is_wysiwyg = "true";
defparam \result_r_tmp[11] .power_up = "low";

dffeas \result_r_tmp[15] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[15]~q ),
	.prn(vcc));
defparam \result_r_tmp[15] .is_wysiwyg = "true";
defparam \result_r_tmp[15] .power_up = "low";

dffeas \result_i_tmp[12] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[12]~q ),
	.prn(vcc));
defparam \result_i_tmp[12] .is_wysiwyg = "true";
defparam \result_i_tmp[12] .power_up = "low";

dffeas \result_r_tmp[12] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[12]~q ),
	.prn(vcc));
defparam \result_r_tmp[12] .is_wysiwyg = "true";
defparam \result_r_tmp[12] .power_up = "low";

dffeas \result_i_tmp[13] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[13]~q ),
	.prn(vcc));
defparam \result_i_tmp[13] .is_wysiwyg = "true";
defparam \result_i_tmp[13] .power_up = "low";

dffeas \result_r_tmp[13] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[13]~q ),
	.prn(vcc));
defparam \result_r_tmp[13] .is_wysiwyg = "true";
defparam \result_r_tmp[13] .power_up = "low";

dffeas \result_i_tmp[14] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[14]~q ),
	.prn(vcc));
defparam \result_i_tmp[14] .is_wysiwyg = "true";
defparam \result_i_tmp[14] .power_up = "low";

dffeas \result_r_tmp[14] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[14]~q ),
	.prn(vcc));
defparam \result_r_tmp[14] .is_wysiwyg = "true";
defparam \result_r_tmp[14] .power_up = "low";

dffeas \result_i_tmp[10] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[10]~q ),
	.prn(vcc));
defparam \result_i_tmp[10] .is_wysiwyg = "true";
defparam \result_i_tmp[10] .power_up = "low";

dffeas \result_r_tmp[10] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[10]~q ),
	.prn(vcc));
defparam \result_r_tmp[10] .is_wysiwyg = "true";
defparam \result_r_tmp[10] .power_up = "low";

dffeas \result_i_tmp[9] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[9]~q ),
	.prn(vcc));
defparam \result_i_tmp[9] .is_wysiwyg = "true";
defparam \result_i_tmp[9] .power_up = "low";

dffeas \result_r_tmp[9] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[9]~q ),
	.prn(vcc));
defparam \result_r_tmp[9] .is_wysiwyg = "true";
defparam \result_r_tmp[9] .power_up = "low";

dffeas \result_i_tmp[8] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[8]~q ),
	.prn(vcc));
defparam \result_i_tmp[8] .is_wysiwyg = "true";
defparam \result_i_tmp[8] .power_up = "low";

dffeas \result_r_tmp[8] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[8]~q ),
	.prn(vcc));
defparam \result_r_tmp[8] .is_wysiwyg = "true";
defparam \result_r_tmp[8] .power_up = "low";

dffeas \result_i_tmp[7] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[7]~q ),
	.prn(vcc));
defparam \result_i_tmp[7] .is_wysiwyg = "true";
defparam \result_i_tmp[7] .power_up = "low";

dffeas \result_r_tmp[7] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[7]~q ),
	.prn(vcc));
defparam \result_r_tmp[7] .is_wysiwyg = "true";
defparam \result_r_tmp[7] .power_up = "low";

dffeas \result_i_tmp[6] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[6]~q ),
	.prn(vcc));
defparam \result_i_tmp[6] .is_wysiwyg = "true";
defparam \result_i_tmp[6] .power_up = "low";

dffeas \result_r_tmp[6] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[6]~q ),
	.prn(vcc));
defparam \result_r_tmp[6] .is_wysiwyg = "true";
defparam \result_r_tmp[6] .power_up = "low";

dffeas \result_i_tmp[5] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[5]~q ),
	.prn(vcc));
defparam \result_i_tmp[5] .is_wysiwyg = "true";
defparam \result_i_tmp[5] .power_up = "low";

dffeas \result_r_tmp[5] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[5]~q ),
	.prn(vcc));
defparam \result_r_tmp[5] .is_wysiwyg = "true";
defparam \result_r_tmp[5] .power_up = "low";

dffeas \result_i_tmp[4] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[4]~q ),
	.prn(vcc));
defparam \result_i_tmp[4] .is_wysiwyg = "true";
defparam \result_i_tmp[4] .power_up = "low";

dffeas \result_r_tmp[4] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[4]~q ),
	.prn(vcc));
defparam \result_r_tmp[4] .is_wysiwyg = "true";
defparam \result_r_tmp[4] .power_up = "low";

dffeas \result_i_tmp[3] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[3]~q ),
	.prn(vcc));
defparam \result_i_tmp[3] .is_wysiwyg = "true";
defparam \result_i_tmp[3] .power_up = "low";

dffeas \result_r_tmp[3] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[3]~q ),
	.prn(vcc));
defparam \result_r_tmp[3] .is_wysiwyg = "true";
defparam \result_r_tmp[3] .power_up = "low";

dffeas \result_i_tmp[2] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[2]~q ),
	.prn(vcc));
defparam \result_i_tmp[2] .is_wysiwyg = "true";
defparam \result_i_tmp[2] .power_up = "low";

dffeas \result_r_tmp[2] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[2]~q ),
	.prn(vcc));
defparam \result_r_tmp[2] .is_wysiwyg = "true";
defparam \result_r_tmp[2] .power_up = "low";

dffeas \result_i_tmp[1] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[1]~q ),
	.prn(vcc));
defparam \result_i_tmp[1] .is_wysiwyg = "true";
defparam \result_i_tmp[1] .power_up = "low";

dffeas \result_r_tmp[1] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[1]~q ),
	.prn(vcc));
defparam \result_r_tmp[1] .is_wysiwyg = "true";
defparam \result_r_tmp[1] .power_up = "low";

dffeas \result_i_tmp[0] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[0]~q ),
	.prn(vcc));
defparam \result_i_tmp[0] .is_wysiwyg = "true";
defparam \result_i_tmp[0] .power_up = "low";

dffeas \result_r_tmp[0] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[0]~q ),
	.prn(vcc));
defparam \result_r_tmp[0] .is_wysiwyg = "true";
defparam \result_r_tmp[0] .power_up = "low";

endmodule

module IFFT_apn_fft_mult_cpx_1 (
	c,
	d,
	global_clock_enable,
	iout_sig2_11,
	iout_sig2_15,
	rout_sig2_11,
	rout_sig2_15,
	iout_sig2_12,
	rout_sig2_12,
	iout_sig2_13,
	rout_sig2_13,
	iout_sig2_14,
	rout_sig2_14,
	iout_sig2_10,
	rout_sig2_10,
	iout_sig2_9,
	rout_sig2_9,
	iout_sig2_8,
	rout_sig2_8,
	b,
	a,
	iout_sig2_7,
	rout_sig2_7,
	iout_sig2_6,
	rout_sig2_6,
	iout_sig2_5,
	rout_sig2_5,
	iout_sig2_4,
	rout_sig2_4,
	iout_sig2_3,
	rout_sig2_3,
	iout_sig2_2,
	rout_sig2_2,
	iout_sig2_1,
	rout_sig2_1,
	iout_sig2_0,
	rout_sig2_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[7:0] c;
input 	[7:0] d;
input 	global_clock_enable;
output 	iout_sig2_11;
output 	iout_sig2_15;
output 	rout_sig2_11;
output 	rout_sig2_15;
output 	iout_sig2_12;
output 	rout_sig2_12;
output 	iout_sig2_13;
output 	rout_sig2_13;
output 	iout_sig2_14;
output 	rout_sig2_14;
output 	iout_sig2_10;
output 	rout_sig2_10;
output 	iout_sig2_9;
output 	rout_sig2_9;
output 	iout_sig2_8;
output 	rout_sig2_8;
input 	[7:0] b;
input 	[7:0] a;
output 	iout_sig2_7;
output 	rout_sig2_7;
output 	iout_sig2_6;
output 	rout_sig2_6;
output 	iout_sig2_5;
output 	rout_sig2_5;
output 	iout_sig2_4;
output 	rout_sig2_4;
output 	iout_sig2_3;
output 	rout_sig2_3;
output 	iout_sig2_2;
output 	rout_sig2_2;
output 	iout_sig2_1;
output 	rout_sig2_1;
output 	iout_sig2_0;
output 	rout_sig2_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~24 ;
wire \Add1~25 ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~28 ;
wire \Add1~29 ;
wire \Add1~30 ;
wire \Add1~31 ;
wire \Add1~32 ;
wire \Add1~33 ;
wire \Add1~34 ;
wire \Add1~35 ;
wire \Add1~36 ;
wire \Add1~37 ;
wire \Add1~38 ;
wire \Add1~39 ;
wire \Add1~40 ;
wire \Add1~41 ;
wire \Add1~42 ;
wire \Add1~43 ;
wire \Add1~44 ;
wire \Add1~45 ;
wire \Add1~46 ;
wire \Add1~47 ;
wire \Add1~48 ;
wire \Add1~49 ;
wire \Add1~50 ;
wire \Add1~51 ;
wire \Add1~52 ;
wire \Add1~53 ;
wire \Add1~54 ;
wire \Add1~55 ;
wire \Add1~56 ;
wire \Add1~57 ;
wire \Add1~58 ;
wire \Add1~59 ;
wire \Add1~60 ;
wire \Add1~61 ;
wire \Add1~62 ;
wire \Add1~63 ;
wire \Add1~64 ;
wire \Add1~65 ;
wire \Add1~66 ;
wire \Add1~67 ;
wire \Add1~68 ;
wire \Add1~69 ;
wire \Add1~70 ;
wire \Add1~71 ;
wire \Add0~24 ;
wire \Add0~25 ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~28 ;
wire \Add0~29 ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~32 ;
wire \Add0~33 ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~36 ;
wire \Add0~37 ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~40 ;
wire \Add0~41 ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~44 ;
wire \Add0~45 ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~48 ;
wire \Add0~49 ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~52 ;
wire \Add0~53 ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~56 ;
wire \Add0~57 ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~60 ;
wire \Add0~61 ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~64 ;
wire \Add0~65 ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~68 ;
wire \Add0~69 ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \c_reg[0]~q ;
wire \c_reg[1]~q ;
wire \c_reg[2]~q ;
wire \c_reg[3]~q ;
wire \c_reg[4]~q ;
wire \c_reg[5]~q ;
wire \c_reg[6]~q ;
wire \c_reg[7]~q ;
wire \b_reg[0]~q ;
wire \b_reg[1]~q ;
wire \b_reg[2]~q ;
wire \b_reg[3]~q ;
wire \b_reg[4]~q ;
wire \b_reg[5]~q ;
wire \b_reg[6]~q ;
wire \b_reg[7]~q ;
wire \d_reg[0]~q ;
wire \d_reg[1]~q ;
wire \d_reg[2]~q ;
wire \d_reg[3]~q ;
wire \d_reg[4]~q ;
wire \d_reg[5]~q ;
wire \d_reg[6]~q ;
wire \d_reg[7]~q ;
wire \a_reg[0]~q ;
wire \a_reg[1]~q ;
wire \a_reg[2]~q ;
wire \a_reg[3]~q ;
wire \a_reg[4]~q ;
wire \a_reg[5]~q ;
wire \a_reg[6]~q ;
wire \a_reg[7]~q ;
wire \Add1~19 ;
wire \iout_sig[11]~q ;
wire \Add1~23 ;
wire \iout_sig[15]~q ;
wire \Add0~19 ;
wire \rout_sig[11]~q ;
wire \Add0~23 ;
wire \rout_sig[15]~q ;
wire \Add1~20 ;
wire \iout_sig[12]~q ;
wire \Add0~20 ;
wire \rout_sig[12]~q ;
wire \Add1~21 ;
wire \iout_sig[13]~q ;
wire \Add0~21 ;
wire \rout_sig[13]~q ;
wire \Add1~22 ;
wire \iout_sig[14]~q ;
wire \Add0~22 ;
wire \rout_sig[14]~q ;
wire \Add1~18 ;
wire \iout_sig[10]~q ;
wire \Add0~18 ;
wire \rout_sig[10]~q ;
wire \Add1~17 ;
wire \iout_sig[9]~q ;
wire \Add0~17 ;
wire \rout_sig[9]~q ;
wire \Add1~16 ;
wire \iout_sig[8]~q ;
wire \Add0~16 ;
wire \rout_sig[8]~q ;
wire \Add1~15 ;
wire \iout_sig[7]~q ;
wire \Add0~15 ;
wire \rout_sig[7]~q ;
wire \Add1~14 ;
wire \iout_sig[6]~q ;
wire \Add0~14 ;
wire \rout_sig[6]~q ;
wire \Add1~13 ;
wire \iout_sig[5]~q ;
wire \Add0~13 ;
wire \rout_sig[5]~q ;
wire \Add1~12 ;
wire \iout_sig[4]~q ;
wire \Add0~12 ;
wire \rout_sig[4]~q ;
wire \Add1~11 ;
wire \iout_sig[3]~q ;
wire \Add0~11 ;
wire \rout_sig[3]~q ;
wire \Add1~10 ;
wire \iout_sig[2]~q ;
wire \Add0~10 ;
wire \rout_sig[2]~q ;
wire \Add1~9 ;
wire \iout_sig[1]~q ;
wire \Add0~9 ;
wire \rout_sig[1]~q ;
wire \Add1~8_resulta ;
wire \iout_sig[0]~q ;
wire \Add0~8_resulta ;
wire \rout_sig[0]~q ;

wire [63:0] \Add1~8_RESULTA_bus ;
wire [63:0] \Add0~8_RESULTA_bus ;

assign \Add1~8_resulta  = \Add1~8_RESULTA_bus [0];
assign \Add1~9  = \Add1~8_RESULTA_bus [1];
assign \Add1~10  = \Add1~8_RESULTA_bus [2];
assign \Add1~11  = \Add1~8_RESULTA_bus [3];
assign \Add1~12  = \Add1~8_RESULTA_bus [4];
assign \Add1~13  = \Add1~8_RESULTA_bus [5];
assign \Add1~14  = \Add1~8_RESULTA_bus [6];
assign \Add1~15  = \Add1~8_RESULTA_bus [7];
assign \Add1~16  = \Add1~8_RESULTA_bus [8];
assign \Add1~17  = \Add1~8_RESULTA_bus [9];
assign \Add1~18  = \Add1~8_RESULTA_bus [10];
assign \Add1~19  = \Add1~8_RESULTA_bus [11];
assign \Add1~20  = \Add1~8_RESULTA_bus [12];
assign \Add1~21  = \Add1~8_RESULTA_bus [13];
assign \Add1~22  = \Add1~8_RESULTA_bus [14];
assign \Add1~23  = \Add1~8_RESULTA_bus [15];
assign \Add1~24  = \Add1~8_RESULTA_bus [16];
assign \Add1~25  = \Add1~8_RESULTA_bus [17];
assign \Add1~26  = \Add1~8_RESULTA_bus [18];
assign \Add1~27  = \Add1~8_RESULTA_bus [19];
assign \Add1~28  = \Add1~8_RESULTA_bus [20];
assign \Add1~29  = \Add1~8_RESULTA_bus [21];
assign \Add1~30  = \Add1~8_RESULTA_bus [22];
assign \Add1~31  = \Add1~8_RESULTA_bus [23];
assign \Add1~32  = \Add1~8_RESULTA_bus [24];
assign \Add1~33  = \Add1~8_RESULTA_bus [25];
assign \Add1~34  = \Add1~8_RESULTA_bus [26];
assign \Add1~35  = \Add1~8_RESULTA_bus [27];
assign \Add1~36  = \Add1~8_RESULTA_bus [28];
assign \Add1~37  = \Add1~8_RESULTA_bus [29];
assign \Add1~38  = \Add1~8_RESULTA_bus [30];
assign \Add1~39  = \Add1~8_RESULTA_bus [31];
assign \Add1~40  = \Add1~8_RESULTA_bus [32];
assign \Add1~41  = \Add1~8_RESULTA_bus [33];
assign \Add1~42  = \Add1~8_RESULTA_bus [34];
assign \Add1~43  = \Add1~8_RESULTA_bus [35];
assign \Add1~44  = \Add1~8_RESULTA_bus [36];
assign \Add1~45  = \Add1~8_RESULTA_bus [37];
assign \Add1~46  = \Add1~8_RESULTA_bus [38];
assign \Add1~47  = \Add1~8_RESULTA_bus [39];
assign \Add1~48  = \Add1~8_RESULTA_bus [40];
assign \Add1~49  = \Add1~8_RESULTA_bus [41];
assign \Add1~50  = \Add1~8_RESULTA_bus [42];
assign \Add1~51  = \Add1~8_RESULTA_bus [43];
assign \Add1~52  = \Add1~8_RESULTA_bus [44];
assign \Add1~53  = \Add1~8_RESULTA_bus [45];
assign \Add1~54  = \Add1~8_RESULTA_bus [46];
assign \Add1~55  = \Add1~8_RESULTA_bus [47];
assign \Add1~56  = \Add1~8_RESULTA_bus [48];
assign \Add1~57  = \Add1~8_RESULTA_bus [49];
assign \Add1~58  = \Add1~8_RESULTA_bus [50];
assign \Add1~59  = \Add1~8_RESULTA_bus [51];
assign \Add1~60  = \Add1~8_RESULTA_bus [52];
assign \Add1~61  = \Add1~8_RESULTA_bus [53];
assign \Add1~62  = \Add1~8_RESULTA_bus [54];
assign \Add1~63  = \Add1~8_RESULTA_bus [55];
assign \Add1~64  = \Add1~8_RESULTA_bus [56];
assign \Add1~65  = \Add1~8_RESULTA_bus [57];
assign \Add1~66  = \Add1~8_RESULTA_bus [58];
assign \Add1~67  = \Add1~8_RESULTA_bus [59];
assign \Add1~68  = \Add1~8_RESULTA_bus [60];
assign \Add1~69  = \Add1~8_RESULTA_bus [61];
assign \Add1~70  = \Add1~8_RESULTA_bus [62];
assign \Add1~71  = \Add1~8_RESULTA_bus [63];

assign \Add0~8_resulta  = \Add0~8_RESULTA_bus [0];
assign \Add0~9  = \Add0~8_RESULTA_bus [1];
assign \Add0~10  = \Add0~8_RESULTA_bus [2];
assign \Add0~11  = \Add0~8_RESULTA_bus [3];
assign \Add0~12  = \Add0~8_RESULTA_bus [4];
assign \Add0~13  = \Add0~8_RESULTA_bus [5];
assign \Add0~14  = \Add0~8_RESULTA_bus [6];
assign \Add0~15  = \Add0~8_RESULTA_bus [7];
assign \Add0~16  = \Add0~8_RESULTA_bus [8];
assign \Add0~17  = \Add0~8_RESULTA_bus [9];
assign \Add0~18  = \Add0~8_RESULTA_bus [10];
assign \Add0~19  = \Add0~8_RESULTA_bus [11];
assign \Add0~20  = \Add0~8_RESULTA_bus [12];
assign \Add0~21  = \Add0~8_RESULTA_bus [13];
assign \Add0~22  = \Add0~8_RESULTA_bus [14];
assign \Add0~23  = \Add0~8_RESULTA_bus [15];
assign \Add0~24  = \Add0~8_RESULTA_bus [16];
assign \Add0~25  = \Add0~8_RESULTA_bus [17];
assign \Add0~26  = \Add0~8_RESULTA_bus [18];
assign \Add0~27  = \Add0~8_RESULTA_bus [19];
assign \Add0~28  = \Add0~8_RESULTA_bus [20];
assign \Add0~29  = \Add0~8_RESULTA_bus [21];
assign \Add0~30  = \Add0~8_RESULTA_bus [22];
assign \Add0~31  = \Add0~8_RESULTA_bus [23];
assign \Add0~32  = \Add0~8_RESULTA_bus [24];
assign \Add0~33  = \Add0~8_RESULTA_bus [25];
assign \Add0~34  = \Add0~8_RESULTA_bus [26];
assign \Add0~35  = \Add0~8_RESULTA_bus [27];
assign \Add0~36  = \Add0~8_RESULTA_bus [28];
assign \Add0~37  = \Add0~8_RESULTA_bus [29];
assign \Add0~38  = \Add0~8_RESULTA_bus [30];
assign \Add0~39  = \Add0~8_RESULTA_bus [31];
assign \Add0~40  = \Add0~8_RESULTA_bus [32];
assign \Add0~41  = \Add0~8_RESULTA_bus [33];
assign \Add0~42  = \Add0~8_RESULTA_bus [34];
assign \Add0~43  = \Add0~8_RESULTA_bus [35];
assign \Add0~44  = \Add0~8_RESULTA_bus [36];
assign \Add0~45  = \Add0~8_RESULTA_bus [37];
assign \Add0~46  = \Add0~8_RESULTA_bus [38];
assign \Add0~47  = \Add0~8_RESULTA_bus [39];
assign \Add0~48  = \Add0~8_RESULTA_bus [40];
assign \Add0~49  = \Add0~8_RESULTA_bus [41];
assign \Add0~50  = \Add0~8_RESULTA_bus [42];
assign \Add0~51  = \Add0~8_RESULTA_bus [43];
assign \Add0~52  = \Add0~8_RESULTA_bus [44];
assign \Add0~53  = \Add0~8_RESULTA_bus [45];
assign \Add0~54  = \Add0~8_RESULTA_bus [46];
assign \Add0~55  = \Add0~8_RESULTA_bus [47];
assign \Add0~56  = \Add0~8_RESULTA_bus [48];
assign \Add0~57  = \Add0~8_RESULTA_bus [49];
assign \Add0~58  = \Add0~8_RESULTA_bus [50];
assign \Add0~59  = \Add0~8_RESULTA_bus [51];
assign \Add0~60  = \Add0~8_RESULTA_bus [52];
assign \Add0~61  = \Add0~8_RESULTA_bus [53];
assign \Add0~62  = \Add0~8_RESULTA_bus [54];
assign \Add0~63  = \Add0~8_RESULTA_bus [55];
assign \Add0~64  = \Add0~8_RESULTA_bus [56];
assign \Add0~65  = \Add0~8_RESULTA_bus [57];
assign \Add0~66  = \Add0~8_RESULTA_bus [58];
assign \Add0~67  = \Add0~8_RESULTA_bus [59];
assign \Add0~68  = \Add0~8_RESULTA_bus [60];
assign \Add0~69  = \Add0~8_RESULTA_bus [61];
assign \Add0~70  = \Add0~8_RESULTA_bus [62];
assign \Add0~71  = \Add0~8_RESULTA_bus [63];

dffeas \iout_sig2[11] (
	.clk(clk),
	.d(\iout_sig[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_11),
	.prn(vcc));
defparam \iout_sig2[11] .is_wysiwyg = "true";
defparam \iout_sig2[11] .power_up = "low";

dffeas \iout_sig2[15] (
	.clk(clk),
	.d(\iout_sig[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_15),
	.prn(vcc));
defparam \iout_sig2[15] .is_wysiwyg = "true";
defparam \iout_sig2[15] .power_up = "low";

dffeas \rout_sig2[11] (
	.clk(clk),
	.d(\rout_sig[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_11),
	.prn(vcc));
defparam \rout_sig2[11] .is_wysiwyg = "true";
defparam \rout_sig2[11] .power_up = "low";

dffeas \rout_sig2[15] (
	.clk(clk),
	.d(\rout_sig[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_15),
	.prn(vcc));
defparam \rout_sig2[15] .is_wysiwyg = "true";
defparam \rout_sig2[15] .power_up = "low";

dffeas \iout_sig2[12] (
	.clk(clk),
	.d(\iout_sig[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_12),
	.prn(vcc));
defparam \iout_sig2[12] .is_wysiwyg = "true";
defparam \iout_sig2[12] .power_up = "low";

dffeas \rout_sig2[12] (
	.clk(clk),
	.d(\rout_sig[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_12),
	.prn(vcc));
defparam \rout_sig2[12] .is_wysiwyg = "true";
defparam \rout_sig2[12] .power_up = "low";

dffeas \iout_sig2[13] (
	.clk(clk),
	.d(\iout_sig[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_13),
	.prn(vcc));
defparam \iout_sig2[13] .is_wysiwyg = "true";
defparam \iout_sig2[13] .power_up = "low";

dffeas \rout_sig2[13] (
	.clk(clk),
	.d(\rout_sig[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_13),
	.prn(vcc));
defparam \rout_sig2[13] .is_wysiwyg = "true";
defparam \rout_sig2[13] .power_up = "low";

dffeas \iout_sig2[14] (
	.clk(clk),
	.d(\iout_sig[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_14),
	.prn(vcc));
defparam \iout_sig2[14] .is_wysiwyg = "true";
defparam \iout_sig2[14] .power_up = "low";

dffeas \rout_sig2[14] (
	.clk(clk),
	.d(\rout_sig[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_14),
	.prn(vcc));
defparam \rout_sig2[14] .is_wysiwyg = "true";
defparam \rout_sig2[14] .power_up = "low";

dffeas \iout_sig2[10] (
	.clk(clk),
	.d(\iout_sig[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_10),
	.prn(vcc));
defparam \iout_sig2[10] .is_wysiwyg = "true";
defparam \iout_sig2[10] .power_up = "low";

dffeas \rout_sig2[10] (
	.clk(clk),
	.d(\rout_sig[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_10),
	.prn(vcc));
defparam \rout_sig2[10] .is_wysiwyg = "true";
defparam \rout_sig2[10] .power_up = "low";

dffeas \iout_sig2[9] (
	.clk(clk),
	.d(\iout_sig[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_9),
	.prn(vcc));
defparam \iout_sig2[9] .is_wysiwyg = "true";
defparam \iout_sig2[9] .power_up = "low";

dffeas \rout_sig2[9] (
	.clk(clk),
	.d(\rout_sig[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_9),
	.prn(vcc));
defparam \rout_sig2[9] .is_wysiwyg = "true";
defparam \rout_sig2[9] .power_up = "low";

dffeas \iout_sig2[8] (
	.clk(clk),
	.d(\iout_sig[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_8),
	.prn(vcc));
defparam \iout_sig2[8] .is_wysiwyg = "true";
defparam \iout_sig2[8] .power_up = "low";

dffeas \rout_sig2[8] (
	.clk(clk),
	.d(\rout_sig[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_8),
	.prn(vcc));
defparam \rout_sig2[8] .is_wysiwyg = "true";
defparam \rout_sig2[8] .power_up = "low";

dffeas \iout_sig2[7] (
	.clk(clk),
	.d(\iout_sig[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_7),
	.prn(vcc));
defparam \iout_sig2[7] .is_wysiwyg = "true";
defparam \iout_sig2[7] .power_up = "low";

dffeas \rout_sig2[7] (
	.clk(clk),
	.d(\rout_sig[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_7),
	.prn(vcc));
defparam \rout_sig2[7] .is_wysiwyg = "true";
defparam \rout_sig2[7] .power_up = "low";

dffeas \iout_sig2[6] (
	.clk(clk),
	.d(\iout_sig[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_6),
	.prn(vcc));
defparam \iout_sig2[6] .is_wysiwyg = "true";
defparam \iout_sig2[6] .power_up = "low";

dffeas \rout_sig2[6] (
	.clk(clk),
	.d(\rout_sig[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_6),
	.prn(vcc));
defparam \rout_sig2[6] .is_wysiwyg = "true";
defparam \rout_sig2[6] .power_up = "low";

dffeas \iout_sig2[5] (
	.clk(clk),
	.d(\iout_sig[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_5),
	.prn(vcc));
defparam \iout_sig2[5] .is_wysiwyg = "true";
defparam \iout_sig2[5] .power_up = "low";

dffeas \rout_sig2[5] (
	.clk(clk),
	.d(\rout_sig[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_5),
	.prn(vcc));
defparam \rout_sig2[5] .is_wysiwyg = "true";
defparam \rout_sig2[5] .power_up = "low";

dffeas \iout_sig2[4] (
	.clk(clk),
	.d(\iout_sig[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_4),
	.prn(vcc));
defparam \iout_sig2[4] .is_wysiwyg = "true";
defparam \iout_sig2[4] .power_up = "low";

dffeas \rout_sig2[4] (
	.clk(clk),
	.d(\rout_sig[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_4),
	.prn(vcc));
defparam \rout_sig2[4] .is_wysiwyg = "true";
defparam \rout_sig2[4] .power_up = "low";

dffeas \iout_sig2[3] (
	.clk(clk),
	.d(\iout_sig[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_3),
	.prn(vcc));
defparam \iout_sig2[3] .is_wysiwyg = "true";
defparam \iout_sig2[3] .power_up = "low";

dffeas \rout_sig2[3] (
	.clk(clk),
	.d(\rout_sig[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_3),
	.prn(vcc));
defparam \rout_sig2[3] .is_wysiwyg = "true";
defparam \rout_sig2[3] .power_up = "low";

dffeas \iout_sig2[2] (
	.clk(clk),
	.d(\iout_sig[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_2),
	.prn(vcc));
defparam \iout_sig2[2] .is_wysiwyg = "true";
defparam \iout_sig2[2] .power_up = "low";

dffeas \rout_sig2[2] (
	.clk(clk),
	.d(\rout_sig[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_2),
	.prn(vcc));
defparam \rout_sig2[2] .is_wysiwyg = "true";
defparam \rout_sig2[2] .power_up = "low";

dffeas \iout_sig2[1] (
	.clk(clk),
	.d(\iout_sig[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_1),
	.prn(vcc));
defparam \iout_sig2[1] .is_wysiwyg = "true";
defparam \iout_sig2[1] .power_up = "low";

dffeas \rout_sig2[1] (
	.clk(clk),
	.d(\rout_sig[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_1),
	.prn(vcc));
defparam \rout_sig2[1] .is_wysiwyg = "true";
defparam \rout_sig2[1] .power_up = "low";

dffeas \iout_sig2[0] (
	.clk(clk),
	.d(\iout_sig[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_0),
	.prn(vcc));
defparam \iout_sig2[0] .is_wysiwyg = "true";
defparam \iout_sig2[0] .power_up = "low";

dffeas \rout_sig2[0] (
	.clk(clk),
	.d(\rout_sig[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_0),
	.prn(vcc));
defparam \rout_sig2[0] .is_wysiwyg = "true";
defparam \rout_sig2[0] .power_up = "low";

dffeas \c_reg[0] (
	.clk(clk),
	.d(c[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[0]~q ),
	.prn(vcc));
defparam \c_reg[0] .is_wysiwyg = "true";
defparam \c_reg[0] .power_up = "low";

dffeas \c_reg[1] (
	.clk(clk),
	.d(c[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[1]~q ),
	.prn(vcc));
defparam \c_reg[1] .is_wysiwyg = "true";
defparam \c_reg[1] .power_up = "low";

dffeas \c_reg[2] (
	.clk(clk),
	.d(c[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[2]~q ),
	.prn(vcc));
defparam \c_reg[2] .is_wysiwyg = "true";
defparam \c_reg[2] .power_up = "low";

dffeas \c_reg[3] (
	.clk(clk),
	.d(c[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[3]~q ),
	.prn(vcc));
defparam \c_reg[3] .is_wysiwyg = "true";
defparam \c_reg[3] .power_up = "low";

dffeas \c_reg[4] (
	.clk(clk),
	.d(c[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[4]~q ),
	.prn(vcc));
defparam \c_reg[4] .is_wysiwyg = "true";
defparam \c_reg[4] .power_up = "low";

dffeas \c_reg[5] (
	.clk(clk),
	.d(c[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[5]~q ),
	.prn(vcc));
defparam \c_reg[5] .is_wysiwyg = "true";
defparam \c_reg[5] .power_up = "low";

dffeas \c_reg[6] (
	.clk(clk),
	.d(c[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[6]~q ),
	.prn(vcc));
defparam \c_reg[6] .is_wysiwyg = "true";
defparam \c_reg[6] .power_up = "low";

dffeas \c_reg[7] (
	.clk(clk),
	.d(c[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[7]~q ),
	.prn(vcc));
defparam \c_reg[7] .is_wysiwyg = "true";
defparam \c_reg[7] .power_up = "low";

dffeas \b_reg[0] (
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[0]~q ),
	.prn(vcc));
defparam \b_reg[0] .is_wysiwyg = "true";
defparam \b_reg[0] .power_up = "low";

dffeas \b_reg[1] (
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[1]~q ),
	.prn(vcc));
defparam \b_reg[1] .is_wysiwyg = "true";
defparam \b_reg[1] .power_up = "low";

dffeas \b_reg[2] (
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[2]~q ),
	.prn(vcc));
defparam \b_reg[2] .is_wysiwyg = "true";
defparam \b_reg[2] .power_up = "low";

dffeas \b_reg[3] (
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[3]~q ),
	.prn(vcc));
defparam \b_reg[3] .is_wysiwyg = "true";
defparam \b_reg[3] .power_up = "low";

dffeas \b_reg[4] (
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[4]~q ),
	.prn(vcc));
defparam \b_reg[4] .is_wysiwyg = "true";
defparam \b_reg[4] .power_up = "low";

dffeas \b_reg[5] (
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[5]~q ),
	.prn(vcc));
defparam \b_reg[5] .is_wysiwyg = "true";
defparam \b_reg[5] .power_up = "low";

dffeas \b_reg[6] (
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[6]~q ),
	.prn(vcc));
defparam \b_reg[6] .is_wysiwyg = "true";
defparam \b_reg[6] .power_up = "low";

dffeas \b_reg[7] (
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[7]~q ),
	.prn(vcc));
defparam \b_reg[7] .is_wysiwyg = "true";
defparam \b_reg[7] .power_up = "low";

dffeas \d_reg[0] (
	.clk(clk),
	.d(d[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[0]~q ),
	.prn(vcc));
defparam \d_reg[0] .is_wysiwyg = "true";
defparam \d_reg[0] .power_up = "low";

dffeas \d_reg[1] (
	.clk(clk),
	.d(d[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[1]~q ),
	.prn(vcc));
defparam \d_reg[1] .is_wysiwyg = "true";
defparam \d_reg[1] .power_up = "low";

dffeas \d_reg[2] (
	.clk(clk),
	.d(d[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[2]~q ),
	.prn(vcc));
defparam \d_reg[2] .is_wysiwyg = "true";
defparam \d_reg[2] .power_up = "low";

dffeas \d_reg[3] (
	.clk(clk),
	.d(d[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[3]~q ),
	.prn(vcc));
defparam \d_reg[3] .is_wysiwyg = "true";
defparam \d_reg[3] .power_up = "low";

dffeas \d_reg[4] (
	.clk(clk),
	.d(d[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[4]~q ),
	.prn(vcc));
defparam \d_reg[4] .is_wysiwyg = "true";
defparam \d_reg[4] .power_up = "low";

dffeas \d_reg[5] (
	.clk(clk),
	.d(d[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[5]~q ),
	.prn(vcc));
defparam \d_reg[5] .is_wysiwyg = "true";
defparam \d_reg[5] .power_up = "low";

dffeas \d_reg[6] (
	.clk(clk),
	.d(d[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[6]~q ),
	.prn(vcc));
defparam \d_reg[6] .is_wysiwyg = "true";
defparam \d_reg[6] .power_up = "low";

dffeas \d_reg[7] (
	.clk(clk),
	.d(d[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[7]~q ),
	.prn(vcc));
defparam \d_reg[7] .is_wysiwyg = "true";
defparam \d_reg[7] .power_up = "low";

dffeas \a_reg[0] (
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[0]~q ),
	.prn(vcc));
defparam \a_reg[0] .is_wysiwyg = "true";
defparam \a_reg[0] .power_up = "low";

dffeas \a_reg[1] (
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[1]~q ),
	.prn(vcc));
defparam \a_reg[1] .is_wysiwyg = "true";
defparam \a_reg[1] .power_up = "low";

dffeas \a_reg[2] (
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[2]~q ),
	.prn(vcc));
defparam \a_reg[2] .is_wysiwyg = "true";
defparam \a_reg[2] .power_up = "low";

dffeas \a_reg[3] (
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[3]~q ),
	.prn(vcc));
defparam \a_reg[3] .is_wysiwyg = "true";
defparam \a_reg[3] .power_up = "low";

dffeas \a_reg[4] (
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[4]~q ),
	.prn(vcc));
defparam \a_reg[4] .is_wysiwyg = "true";
defparam \a_reg[4] .power_up = "low";

dffeas \a_reg[5] (
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[5]~q ),
	.prn(vcc));
defparam \a_reg[5] .is_wysiwyg = "true";
defparam \a_reg[5] .power_up = "low";

dffeas \a_reg[6] (
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[6]~q ),
	.prn(vcc));
defparam \a_reg[6] .is_wysiwyg = "true";
defparam \a_reg[6] .power_up = "low";

dffeas \a_reg[7] (
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[7]~q ),
	.prn(vcc));
defparam \a_reg[7] .is_wysiwyg = "true";
defparam \a_reg[7] .power_up = "low";

cyclonev_mac \Add1~8 (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\c_reg[7]~q ,\c_reg[6]~q ,\c_reg[5]~q ,\c_reg[4]~q ,\c_reg[3]~q ,\c_reg[2]~q ,\c_reg[1]~q ,\c_reg[0]~q }),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\b_reg[7]~q ,\b_reg[6]~q ,\b_reg[5]~q ,\b_reg[4]~q ,\b_reg[3]~q ,\b_reg[2]~q ,\b_reg[1]~q ,\b_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_reg[7]~q ,\d_reg[6]~q ,\d_reg[5]~q ,\d_reg[4]~q ,\d_reg[3]~q ,\d_reg[2]~q ,\d_reg[1]~q ,\d_reg[0]~q }),
	.by({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\a_reg[7]~q ,\a_reg[6]~q ,\a_reg[5]~q ,\a_reg[4]~q ,\a_reg[3]~q ,\a_reg[2]~q ,\a_reg[1]~q ,\a_reg[0]~q }),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Add1~8_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Add1~8 .accumulate_clock = "none";
defparam \Add1~8 .ax_clock = "none";
defparam \Add1~8 .ax_width = 8;
defparam \Add1~8 .ay_scan_in_clock = "none";
defparam \Add1~8 .ay_scan_in_width = 8;
defparam \Add1~8 .ay_use_scan_in = "false";
defparam \Add1~8 .az_clock = "none";
defparam \Add1~8 .bx_clock = "none";
defparam \Add1~8 .bx_width = 8;
defparam \Add1~8 .by_clock = "none";
defparam \Add1~8 .by_use_scan_in = "false";
defparam \Add1~8 .by_width = 8;
defparam \Add1~8 .bz_clock = "none";
defparam \Add1~8 .coef_a_0 = 0;
defparam \Add1~8 .coef_a_1 = 0;
defparam \Add1~8 .coef_a_2 = 0;
defparam \Add1~8 .coef_a_3 = 0;
defparam \Add1~8 .coef_a_4 = 0;
defparam \Add1~8 .coef_a_5 = 0;
defparam \Add1~8 .coef_a_6 = 0;
defparam \Add1~8 .coef_a_7 = 0;
defparam \Add1~8 .coef_b_0 = 0;
defparam \Add1~8 .coef_b_1 = 0;
defparam \Add1~8 .coef_b_2 = 0;
defparam \Add1~8 .coef_b_3 = 0;
defparam \Add1~8 .coef_b_4 = 0;
defparam \Add1~8 .coef_b_5 = 0;
defparam \Add1~8 .coef_b_6 = 0;
defparam \Add1~8 .coef_b_7 = 0;
defparam \Add1~8 .coef_sel_a_clock = "none";
defparam \Add1~8 .coef_sel_b_clock = "none";
defparam \Add1~8 .delay_scan_out_ay = "false";
defparam \Add1~8 .delay_scan_out_by = "false";
defparam \Add1~8 .enable_double_accum = "false";
defparam \Add1~8 .load_const_clock = "none";
defparam \Add1~8 .load_const_value = 0;
defparam \Add1~8 .mode_sub_location = 0;
defparam \Add1~8 .negate_clock = "none";
defparam \Add1~8 .operand_source_max = "input";
defparam \Add1~8 .operand_source_may = "input";
defparam \Add1~8 .operand_source_mbx = "input";
defparam \Add1~8 .operand_source_mby = "input";
defparam \Add1~8 .operation_mode = "m18x18_sumof2";
defparam \Add1~8 .output_clock = "none";
defparam \Add1~8 .preadder_subtract_a = "false";
defparam \Add1~8 .preadder_subtract_b = "false";
defparam \Add1~8 .result_a_width = 64;
defparam \Add1~8 .signed_max = "true";
defparam \Add1~8 .signed_may = "true";
defparam \Add1~8 .signed_mbx = "true";
defparam \Add1~8 .signed_mby = "true";
defparam \Add1~8 .sub_clock = "none";
defparam \Add1~8 .use_chainadder = "false";

dffeas \iout_sig[11] (
	.clk(clk),
	.d(\Add1~19 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[11]~q ),
	.prn(vcc));
defparam \iout_sig[11] .is_wysiwyg = "true";
defparam \iout_sig[11] .power_up = "low";

dffeas \iout_sig[15] (
	.clk(clk),
	.d(\Add1~23 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[15]~q ),
	.prn(vcc));
defparam \iout_sig[15] .is_wysiwyg = "true";
defparam \iout_sig[15] .power_up = "low";

cyclonev_mac \Add0~8 (
	.sub(vcc),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_reg[7]~q ,\d_reg[6]~q ,\d_reg[5]~q ,\d_reg[4]~q ,\d_reg[3]~q ,\d_reg[2]~q ,\d_reg[1]~q ,\d_reg[0]~q }),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\b_reg[7]~q ,\b_reg[6]~q ,\b_reg[5]~q ,\b_reg[4]~q ,\b_reg[3]~q ,\b_reg[2]~q ,\b_reg[1]~q ,\b_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\c_reg[7]~q ,\c_reg[6]~q ,\c_reg[5]~q ,\c_reg[4]~q ,\c_reg[3]~q ,\c_reg[2]~q ,\c_reg[1]~q ,\c_reg[0]~q }),
	.by({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\a_reg[7]~q ,\a_reg[6]~q ,\a_reg[5]~q ,\a_reg[4]~q ,\a_reg[3]~q ,\a_reg[2]~q ,\a_reg[1]~q ,\a_reg[0]~q }),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Add0~8_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Add0~8 .accumulate_clock = "none";
defparam \Add0~8 .ax_clock = "none";
defparam \Add0~8 .ax_width = 8;
defparam \Add0~8 .ay_scan_in_clock = "none";
defparam \Add0~8 .ay_scan_in_width = 8;
defparam \Add0~8 .ay_use_scan_in = "false";
defparam \Add0~8 .az_clock = "none";
defparam \Add0~8 .bx_clock = "none";
defparam \Add0~8 .bx_width = 8;
defparam \Add0~8 .by_clock = "none";
defparam \Add0~8 .by_use_scan_in = "false";
defparam \Add0~8 .by_width = 8;
defparam \Add0~8 .bz_clock = "none";
defparam \Add0~8 .coef_a_0 = 0;
defparam \Add0~8 .coef_a_1 = 0;
defparam \Add0~8 .coef_a_2 = 0;
defparam \Add0~8 .coef_a_3 = 0;
defparam \Add0~8 .coef_a_4 = 0;
defparam \Add0~8 .coef_a_5 = 0;
defparam \Add0~8 .coef_a_6 = 0;
defparam \Add0~8 .coef_a_7 = 0;
defparam \Add0~8 .coef_b_0 = 0;
defparam \Add0~8 .coef_b_1 = 0;
defparam \Add0~8 .coef_b_2 = 0;
defparam \Add0~8 .coef_b_3 = 0;
defparam \Add0~8 .coef_b_4 = 0;
defparam \Add0~8 .coef_b_5 = 0;
defparam \Add0~8 .coef_b_6 = 0;
defparam \Add0~8 .coef_b_7 = 0;
defparam \Add0~8 .coef_sel_a_clock = "none";
defparam \Add0~8 .coef_sel_b_clock = "none";
defparam \Add0~8 .delay_scan_out_ay = "false";
defparam \Add0~8 .delay_scan_out_by = "false";
defparam \Add0~8 .enable_double_accum = "false";
defparam \Add0~8 .load_const_clock = "none";
defparam \Add0~8 .load_const_value = 0;
defparam \Add0~8 .mode_sub_location = 0;
defparam \Add0~8 .negate_clock = "none";
defparam \Add0~8 .operand_source_max = "input";
defparam \Add0~8 .operand_source_may = "input";
defparam \Add0~8 .operand_source_mbx = "input";
defparam \Add0~8 .operand_source_mby = "input";
defparam \Add0~8 .operation_mode = "m18x18_sumof2";
defparam \Add0~8 .output_clock = "none";
defparam \Add0~8 .preadder_subtract_a = "false";
defparam \Add0~8 .preadder_subtract_b = "false";
defparam \Add0~8 .result_a_width = 64;
defparam \Add0~8 .signed_max = "true";
defparam \Add0~8 .signed_may = "true";
defparam \Add0~8 .signed_mbx = "true";
defparam \Add0~8 .signed_mby = "true";
defparam \Add0~8 .sub_clock = "none";
defparam \Add0~8 .use_chainadder = "false";

dffeas \rout_sig[11] (
	.clk(clk),
	.d(\Add0~19 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[11]~q ),
	.prn(vcc));
defparam \rout_sig[11] .is_wysiwyg = "true";
defparam \rout_sig[11] .power_up = "low";

dffeas \rout_sig[15] (
	.clk(clk),
	.d(\Add0~23 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[15]~q ),
	.prn(vcc));
defparam \rout_sig[15] .is_wysiwyg = "true";
defparam \rout_sig[15] .power_up = "low";

dffeas \iout_sig[12] (
	.clk(clk),
	.d(\Add1~20 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[12]~q ),
	.prn(vcc));
defparam \iout_sig[12] .is_wysiwyg = "true";
defparam \iout_sig[12] .power_up = "low";

dffeas \rout_sig[12] (
	.clk(clk),
	.d(\Add0~20 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[12]~q ),
	.prn(vcc));
defparam \rout_sig[12] .is_wysiwyg = "true";
defparam \rout_sig[12] .power_up = "low";

dffeas \iout_sig[13] (
	.clk(clk),
	.d(\Add1~21 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[13]~q ),
	.prn(vcc));
defparam \iout_sig[13] .is_wysiwyg = "true";
defparam \iout_sig[13] .power_up = "low";

dffeas \rout_sig[13] (
	.clk(clk),
	.d(\Add0~21 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[13]~q ),
	.prn(vcc));
defparam \rout_sig[13] .is_wysiwyg = "true";
defparam \rout_sig[13] .power_up = "low";

dffeas \iout_sig[14] (
	.clk(clk),
	.d(\Add1~22 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[14]~q ),
	.prn(vcc));
defparam \iout_sig[14] .is_wysiwyg = "true";
defparam \iout_sig[14] .power_up = "low";

dffeas \rout_sig[14] (
	.clk(clk),
	.d(\Add0~22 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[14]~q ),
	.prn(vcc));
defparam \rout_sig[14] .is_wysiwyg = "true";
defparam \rout_sig[14] .power_up = "low";

dffeas \iout_sig[10] (
	.clk(clk),
	.d(\Add1~18 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[10]~q ),
	.prn(vcc));
defparam \iout_sig[10] .is_wysiwyg = "true";
defparam \iout_sig[10] .power_up = "low";

dffeas \rout_sig[10] (
	.clk(clk),
	.d(\Add0~18 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[10]~q ),
	.prn(vcc));
defparam \rout_sig[10] .is_wysiwyg = "true";
defparam \rout_sig[10] .power_up = "low";

dffeas \iout_sig[9] (
	.clk(clk),
	.d(\Add1~17 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[9]~q ),
	.prn(vcc));
defparam \iout_sig[9] .is_wysiwyg = "true";
defparam \iout_sig[9] .power_up = "low";

dffeas \rout_sig[9] (
	.clk(clk),
	.d(\Add0~17 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[9]~q ),
	.prn(vcc));
defparam \rout_sig[9] .is_wysiwyg = "true";
defparam \rout_sig[9] .power_up = "low";

dffeas \iout_sig[8] (
	.clk(clk),
	.d(\Add1~16 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[8]~q ),
	.prn(vcc));
defparam \iout_sig[8] .is_wysiwyg = "true";
defparam \iout_sig[8] .power_up = "low";

dffeas \rout_sig[8] (
	.clk(clk),
	.d(\Add0~16 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[8]~q ),
	.prn(vcc));
defparam \rout_sig[8] .is_wysiwyg = "true";
defparam \rout_sig[8] .power_up = "low";

dffeas \iout_sig[7] (
	.clk(clk),
	.d(\Add1~15 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[7]~q ),
	.prn(vcc));
defparam \iout_sig[7] .is_wysiwyg = "true";
defparam \iout_sig[7] .power_up = "low";

dffeas \rout_sig[7] (
	.clk(clk),
	.d(\Add0~15 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[7]~q ),
	.prn(vcc));
defparam \rout_sig[7] .is_wysiwyg = "true";
defparam \rout_sig[7] .power_up = "low";

dffeas \iout_sig[6] (
	.clk(clk),
	.d(\Add1~14 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[6]~q ),
	.prn(vcc));
defparam \iout_sig[6] .is_wysiwyg = "true";
defparam \iout_sig[6] .power_up = "low";

dffeas \rout_sig[6] (
	.clk(clk),
	.d(\Add0~14 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[6]~q ),
	.prn(vcc));
defparam \rout_sig[6] .is_wysiwyg = "true";
defparam \rout_sig[6] .power_up = "low";

dffeas \iout_sig[5] (
	.clk(clk),
	.d(\Add1~13 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[5]~q ),
	.prn(vcc));
defparam \iout_sig[5] .is_wysiwyg = "true";
defparam \iout_sig[5] .power_up = "low";

dffeas \rout_sig[5] (
	.clk(clk),
	.d(\Add0~13 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[5]~q ),
	.prn(vcc));
defparam \rout_sig[5] .is_wysiwyg = "true";
defparam \rout_sig[5] .power_up = "low";

dffeas \iout_sig[4] (
	.clk(clk),
	.d(\Add1~12 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[4]~q ),
	.prn(vcc));
defparam \iout_sig[4] .is_wysiwyg = "true";
defparam \iout_sig[4] .power_up = "low";

dffeas \rout_sig[4] (
	.clk(clk),
	.d(\Add0~12 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[4]~q ),
	.prn(vcc));
defparam \rout_sig[4] .is_wysiwyg = "true";
defparam \rout_sig[4] .power_up = "low";

dffeas \iout_sig[3] (
	.clk(clk),
	.d(\Add1~11 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[3]~q ),
	.prn(vcc));
defparam \iout_sig[3] .is_wysiwyg = "true";
defparam \iout_sig[3] .power_up = "low";

dffeas \rout_sig[3] (
	.clk(clk),
	.d(\Add0~11 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[3]~q ),
	.prn(vcc));
defparam \rout_sig[3] .is_wysiwyg = "true";
defparam \rout_sig[3] .power_up = "low";

dffeas \iout_sig[2] (
	.clk(clk),
	.d(\Add1~10 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[2]~q ),
	.prn(vcc));
defparam \iout_sig[2] .is_wysiwyg = "true";
defparam \iout_sig[2] .power_up = "low";

dffeas \rout_sig[2] (
	.clk(clk),
	.d(\Add0~10 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[2]~q ),
	.prn(vcc));
defparam \rout_sig[2] .is_wysiwyg = "true";
defparam \rout_sig[2] .power_up = "low";

dffeas \iout_sig[1] (
	.clk(clk),
	.d(\Add1~9 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[1]~q ),
	.prn(vcc));
defparam \iout_sig[1] .is_wysiwyg = "true";
defparam \iout_sig[1] .power_up = "low";

dffeas \rout_sig[1] (
	.clk(clk),
	.d(\Add0~9 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[1]~q ),
	.prn(vcc));
defparam \rout_sig[1] .is_wysiwyg = "true";
defparam \rout_sig[1] .power_up = "low";

dffeas \iout_sig[0] (
	.clk(clk),
	.d(\Add1~8_resulta ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[0]~q ),
	.prn(vcc));
defparam \iout_sig[0] .is_wysiwyg = "true";
defparam \iout_sig[0] .power_up = "low";

dffeas \rout_sig[0] (
	.clk(clk),
	.d(\Add0~8_resulta ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[0]~q ),
	.prn(vcc));
defparam \rout_sig[0] .is_wysiwyg = "true";
defparam \rout_sig[0] .power_up = "low";

endmodule

module IFFT_asj_fft_pround_2 (
	global_clock_enable,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_3 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_r_tmp_8(result_r_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_r_tmp_7(result_r_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_3 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_8gj_2 auto_generated(
	.clken(clken),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_r_tmp_8(result_r_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_r_tmp_7(result_r_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.clock(clock));

endmodule

module IFFT_add_sub_8gj_2 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_3 (
	global_clock_enable,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_4 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_i_tmp_8(result_i_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_i_tmp_7(result_i_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_4 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_8gj_3 auto_generated(
	.clken(clken),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_i_tmp_8(result_i_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_i_tmp_7(result_i_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.clock(clock));

endmodule

module IFFT_add_sub_8gj_3 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm2|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl_2 (
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_4_1,
	tdl_arr_5_1,
	tdl_arr_6_1,
	data_in,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_4_1;
output 	tdl_arr_5_1;
output 	tdl_arr_6_1;
input 	[7:0] data_in;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][3]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;


dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_3 (
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_4_1,
	tdl_arr_5_1,
	tdl_arr_6_1,
	data_in,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_4_1;
output 	tdl_arr_5_1;
output 	tdl_arr_6_1;
input 	[7:0] data_in;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][3]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;


dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

endmodule

module IFFT_apn_fft_cmult_cpx2_2 (
	twiddle_data207,
	twiddle_data210,
	twiddle_data211,
	twiddle_data212,
	twiddle_data213,
	twiddle_data214,
	twiddle_data215,
	twiddle_data216,
	twiddle_data217,
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_3_11,
	tdl_arr_7_11,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_5_1,
	tdl_arr_5_11,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_2_1,
	tdl_arr_2_11,
	tdl_arr_1_1,
	tdl_arr_1_11,
	tdl_arr_0_1,
	tdl_arr_0_11,
	twiddle_data200,
	twiddle_data201,
	twiddle_data202,
	twiddle_data203,
	twiddle_data204,
	twiddle_data205,
	twiddle_data206,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	twiddle_data207;
input 	twiddle_data210;
input 	twiddle_data211;
input 	twiddle_data212;
input 	twiddle_data213;
input 	twiddle_data214;
input 	twiddle_data215;
input 	twiddle_data216;
input 	twiddle_data217;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_3_11;
output 	tdl_arr_7_11;
output 	tdl_arr_4_1;
output 	tdl_arr_4_11;
output 	tdl_arr_5_1;
output 	tdl_arr_5_11;
output 	tdl_arr_6_1;
output 	tdl_arr_6_11;
output 	tdl_arr_2_1;
output 	tdl_arr_2_11;
output 	tdl_arr_1_1;
output 	tdl_arr_1_11;
output 	tdl_arr_0_1;
output 	tdl_arr_0_11;
input 	twiddle_data200;
input 	twiddle_data201;
input 	twiddle_data202;
input 	twiddle_data203;
input 	twiddle_data204;
input 	twiddle_data205;
input 	twiddle_data206;
input 	pipeline_dffe_2;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ;
wire \result_i_tmp[11]~q ;
wire \result_i_tmp[15]~q ;
wire \result_r_tmp[11]~q ;
wire \result_r_tmp[15]~q ;
wire \result_i_tmp[12]~q ;
wire \result_r_tmp[12]~q ;
wire \result_i_tmp[13]~q ;
wire \result_r_tmp[13]~q ;
wire \result_i_tmp[14]~q ;
wire \result_r_tmp[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ;
wire \result_i_tmp[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ;
wire \result_r_tmp[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ;
wire \result_i_tmp[9]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ;
wire \result_r_tmp[9]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ;
wire \result_i_tmp[8]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ;
wire \result_r_tmp[8]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ;
wire \result_i_tmp[7]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ;
wire \result_r_tmp[7]~q ;
wire \u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ;
wire \result_i_tmp[6]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ;
wire \result_r_tmp[6]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ;
wire \result_i_tmp[5]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ;
wire \result_r_tmp[5]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ;
wire \result_i_tmp[4]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ;
wire \result_r_tmp[4]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ;
wire \result_i_tmp[3]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ;
wire \result_r_tmp[3]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ;
wire \result_i_tmp[2]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ;
wire \result_r_tmp[2]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ;
wire \result_i_tmp[1]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ;
wire \result_r_tmp[1]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ;
wire \result_i_tmp[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ;
wire \result_r_tmp[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ;
wire \gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ;


IFFT_asj_fft_tdl_4 imag_delay(
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_1),
	.tdl_arr_7_1(tdl_arr_7_1),
	.tdl_arr_4_1(tdl_arr_4_1),
	.tdl_arr_5_1(tdl_arr_5_1),
	.tdl_arr_6_1(tdl_arr_6_1),
	.data_in({\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,
\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ,
\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ,\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q }),
	.tdl_arr_2_1(tdl_arr_2_1),
	.tdl_arr_1_1(tdl_arr_1_1),
	.tdl_arr_0_1(tdl_arr_0_1),
	.clk(clk));

IFFT_asj_fft_tdl_5 real_delay(
	.global_clock_enable(global_clock_enable),
	.tdl_arr_3_1(tdl_arr_3_11),
	.tdl_arr_7_1(tdl_arr_7_11),
	.tdl_arr_4_1(tdl_arr_4_11),
	.tdl_arr_5_1(tdl_arr_5_11),
	.tdl_arr_6_1(tdl_arr_6_11),
	.data_in({\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ,
\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ,
\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ,\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q }),
	.tdl_arr_2_1(tdl_arr_2_11),
	.tdl_arr_1_1(tdl_arr_1_11),
	.tdl_arr_0_1(tdl_arr_0_11),
	.clk(clk));

IFFT_asj_fft_pround_5 u1(
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_11(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_i_tmp_11(\result_i_tmp[11]~q ),
	.result_i_tmp_15(\result_i_tmp[15]~q ),
	.result_i_tmp_12(\result_i_tmp[12]~q ),
	.result_i_tmp_13(\result_i_tmp[13]~q ),
	.result_i_tmp_14(\result_i_tmp[14]~q ),
	.result_i_tmp_10(\result_i_tmp[10]~q ),
	.result_i_tmp_9(\result_i_tmp[9]~q ),
	.pipeline_dffe_10(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.result_i_tmp_8(\result_i_tmp[8]~q ),
	.pipeline_dffe_9(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.result_i_tmp_7(\result_i_tmp[7]~q ),
	.pipeline_dffe_8(\u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.result_i_tmp_6(\result_i_tmp[6]~q ),
	.result_i_tmp_5(\result_i_tmp[5]~q ),
	.result_i_tmp_4(\result_i_tmp[4]~q ),
	.result_i_tmp_3(\result_i_tmp[3]~q ),
	.result_i_tmp_2(\result_i_tmp[2]~q ),
	.result_i_tmp_1(\result_i_tmp[1]~q ),
	.result_i_tmp_0(\result_i_tmp[0]~q ),
	.clk(clk));

IFFT_asj_fft_pround_4 u0(
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_11(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_15(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14]~q ),
	.result_r_tmp_11(\result_r_tmp[11]~q ),
	.result_r_tmp_15(\result_r_tmp[15]~q ),
	.result_r_tmp_12(\result_r_tmp[12]~q ),
	.result_r_tmp_13(\result_r_tmp[13]~q ),
	.result_r_tmp_14(\result_r_tmp[14]~q ),
	.result_r_tmp_10(\result_r_tmp[10]~q ),
	.result_r_tmp_9(\result_r_tmp[9]~q ),
	.pipeline_dffe_10(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10]~q ),
	.result_r_tmp_8(\result_r_tmp[8]~q ),
	.pipeline_dffe_9(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.result_r_tmp_7(\result_r_tmp[7]~q ),
	.pipeline_dffe_8(\u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.result_r_tmp_6(\result_r_tmp[6]~q ),
	.result_r_tmp_5(\result_r_tmp[5]~q ),
	.result_r_tmp_4(\result_r_tmp[4]~q ),
	.result_r_tmp_3(\result_r_tmp[3]~q ),
	.result_r_tmp_2(\result_r_tmp[2]~q ),
	.result_r_tmp_1(\result_r_tmp[1]~q ),
	.result_r_tmp_0(\result_r_tmp[0]~q ),
	.clk(clk));

IFFT_apn_fft_mult_cpx_2 \gen_infr_4cpx:calc_mult_4cpx (
	.c({twiddle_data207,twiddle_data206,twiddle_data205,twiddle_data204,twiddle_data203,twiddle_data202,twiddle_data201,twiddle_data200}),
	.d({twiddle_data217,twiddle_data216,twiddle_data215,twiddle_data214,twiddle_data213,twiddle_data212,twiddle_data211,twiddle_data210}),
	.global_clock_enable(global_clock_enable),
	.iout_sig2_11(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ),
	.iout_sig2_15(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ),
	.rout_sig2_11(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ),
	.rout_sig2_15(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ),
	.iout_sig2_12(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ),
	.rout_sig2_12(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ),
	.iout_sig2_13(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ),
	.rout_sig2_13(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ),
	.iout_sig2_14(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ),
	.rout_sig2_14(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ),
	.iout_sig2_10(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ),
	.rout_sig2_10(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ),
	.iout_sig2_9(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ),
	.rout_sig2_9(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ),
	.iout_sig2_8(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ),
	.rout_sig2_8(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ),
	.b({pipeline_dffe_9,pipeline_dffe_8,pipeline_dffe_7,pipeline_dffe_6,pipeline_dffe_5,pipeline_dffe_4,pipeline_dffe_3,pipeline_dffe_2}),
	.a({pipeline_dffe_91,pipeline_dffe_81,pipeline_dffe_71,pipeline_dffe_61,pipeline_dffe_51,pipeline_dffe_41,pipeline_dffe_31,pipeline_dffe_21}),
	.iout_sig2_7(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ),
	.rout_sig2_7(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ),
	.iout_sig2_6(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ),
	.rout_sig2_6(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ),
	.iout_sig2_5(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ),
	.rout_sig2_5(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ),
	.iout_sig2_4(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ),
	.rout_sig2_4(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ),
	.iout_sig2_3(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ),
	.rout_sig2_3(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ),
	.iout_sig2_2(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ),
	.rout_sig2_2(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ),
	.iout_sig2_1(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ),
	.rout_sig2_1(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ),
	.iout_sig2_0(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ),
	.rout_sig2_0(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ),
	.clk(clk),
	.reset(reset));

dffeas \result_i_tmp[11] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[11]~q ),
	.prn(vcc));
defparam \result_i_tmp[11] .is_wysiwyg = "true";
defparam \result_i_tmp[11] .power_up = "low";

dffeas \result_i_tmp[15] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[15]~q ),
	.prn(vcc));
defparam \result_i_tmp[15] .is_wysiwyg = "true";
defparam \result_i_tmp[15] .power_up = "low";

dffeas \result_r_tmp[11] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[11]~q ),
	.prn(vcc));
defparam \result_r_tmp[11] .is_wysiwyg = "true";
defparam \result_r_tmp[11] .power_up = "low";

dffeas \result_r_tmp[15] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[15]~q ),
	.prn(vcc));
defparam \result_r_tmp[15] .is_wysiwyg = "true";
defparam \result_r_tmp[15] .power_up = "low";

dffeas \result_i_tmp[12] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[12]~q ),
	.prn(vcc));
defparam \result_i_tmp[12] .is_wysiwyg = "true";
defparam \result_i_tmp[12] .power_up = "low";

dffeas \result_r_tmp[12] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[12]~q ),
	.prn(vcc));
defparam \result_r_tmp[12] .is_wysiwyg = "true";
defparam \result_r_tmp[12] .power_up = "low";

dffeas \result_i_tmp[13] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[13]~q ),
	.prn(vcc));
defparam \result_i_tmp[13] .is_wysiwyg = "true";
defparam \result_i_tmp[13] .power_up = "low";

dffeas \result_r_tmp[13] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[13]~q ),
	.prn(vcc));
defparam \result_r_tmp[13] .is_wysiwyg = "true";
defparam \result_r_tmp[13] .power_up = "low";

dffeas \result_i_tmp[14] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[14]~q ),
	.prn(vcc));
defparam \result_i_tmp[14] .is_wysiwyg = "true";
defparam \result_i_tmp[14] .power_up = "low";

dffeas \result_r_tmp[14] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[14]~q ),
	.prn(vcc));
defparam \result_r_tmp[14] .is_wysiwyg = "true";
defparam \result_r_tmp[14] .power_up = "low";

dffeas \result_i_tmp[10] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[10]~q ),
	.prn(vcc));
defparam \result_i_tmp[10] .is_wysiwyg = "true";
defparam \result_i_tmp[10] .power_up = "low";

dffeas \result_r_tmp[10] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[10]~q ),
	.prn(vcc));
defparam \result_r_tmp[10] .is_wysiwyg = "true";
defparam \result_r_tmp[10] .power_up = "low";

dffeas \result_i_tmp[9] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[9]~q ),
	.prn(vcc));
defparam \result_i_tmp[9] .is_wysiwyg = "true";
defparam \result_i_tmp[9] .power_up = "low";

dffeas \result_r_tmp[9] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[9]~q ),
	.prn(vcc));
defparam \result_r_tmp[9] .is_wysiwyg = "true";
defparam \result_r_tmp[9] .power_up = "low";

dffeas \result_i_tmp[8] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[8]~q ),
	.prn(vcc));
defparam \result_i_tmp[8] .is_wysiwyg = "true";
defparam \result_i_tmp[8] .power_up = "low";

dffeas \result_r_tmp[8] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[8]~q ),
	.prn(vcc));
defparam \result_r_tmp[8] .is_wysiwyg = "true";
defparam \result_r_tmp[8] .power_up = "low";

dffeas \result_i_tmp[7] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[7]~q ),
	.prn(vcc));
defparam \result_i_tmp[7] .is_wysiwyg = "true";
defparam \result_i_tmp[7] .power_up = "low";

dffeas \result_r_tmp[7] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[7]~q ),
	.prn(vcc));
defparam \result_r_tmp[7] .is_wysiwyg = "true";
defparam \result_r_tmp[7] .power_up = "low";

dffeas \result_i_tmp[6] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[6]~q ),
	.prn(vcc));
defparam \result_i_tmp[6] .is_wysiwyg = "true";
defparam \result_i_tmp[6] .power_up = "low";

dffeas \result_r_tmp[6] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[6]~q ),
	.prn(vcc));
defparam \result_r_tmp[6] .is_wysiwyg = "true";
defparam \result_r_tmp[6] .power_up = "low";

dffeas \result_i_tmp[5] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[5]~q ),
	.prn(vcc));
defparam \result_i_tmp[5] .is_wysiwyg = "true";
defparam \result_i_tmp[5] .power_up = "low";

dffeas \result_r_tmp[5] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[5]~q ),
	.prn(vcc));
defparam \result_r_tmp[5] .is_wysiwyg = "true";
defparam \result_r_tmp[5] .power_up = "low";

dffeas \result_i_tmp[4] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[4]~q ),
	.prn(vcc));
defparam \result_i_tmp[4] .is_wysiwyg = "true";
defparam \result_i_tmp[4] .power_up = "low";

dffeas \result_r_tmp[4] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[4]~q ),
	.prn(vcc));
defparam \result_r_tmp[4] .is_wysiwyg = "true";
defparam \result_r_tmp[4] .power_up = "low";

dffeas \result_i_tmp[3] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[3]~q ),
	.prn(vcc));
defparam \result_i_tmp[3] .is_wysiwyg = "true";
defparam \result_i_tmp[3] .power_up = "low";

dffeas \result_r_tmp[3] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[3]~q ),
	.prn(vcc));
defparam \result_r_tmp[3] .is_wysiwyg = "true";
defparam \result_r_tmp[3] .power_up = "low";

dffeas \result_i_tmp[2] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[2]~q ),
	.prn(vcc));
defparam \result_i_tmp[2] .is_wysiwyg = "true";
defparam \result_i_tmp[2] .power_up = "low";

dffeas \result_r_tmp[2] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[2]~q ),
	.prn(vcc));
defparam \result_r_tmp[2] .is_wysiwyg = "true";
defparam \result_r_tmp[2] .power_up = "low";

dffeas \result_i_tmp[1] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[1]~q ),
	.prn(vcc));
defparam \result_i_tmp[1] .is_wysiwyg = "true";
defparam \result_i_tmp[1] .power_up = "low";

dffeas \result_r_tmp[1] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[1]~q ),
	.prn(vcc));
defparam \result_r_tmp[1] .is_wysiwyg = "true";
defparam \result_r_tmp[1] .power_up = "low";

dffeas \result_i_tmp[0] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|iout_sig2[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_i_tmp[0]~q ),
	.prn(vcc));
defparam \result_i_tmp[0] .is_wysiwyg = "true";
defparam \result_i_tmp[0] .power_up = "low";

dffeas \result_r_tmp[0] (
	.clk(clk),
	.d(\gen_infr_4cpx:calc_mult_4cpx|rout_sig2[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_r_tmp[0]~q ),
	.prn(vcc));
defparam \result_r_tmp[0] .is_wysiwyg = "true";
defparam \result_r_tmp[0] .power_up = "low";

endmodule

module IFFT_apn_fft_mult_cpx_2 (
	c,
	d,
	global_clock_enable,
	iout_sig2_11,
	iout_sig2_15,
	rout_sig2_11,
	rout_sig2_15,
	iout_sig2_12,
	rout_sig2_12,
	iout_sig2_13,
	rout_sig2_13,
	iout_sig2_14,
	rout_sig2_14,
	iout_sig2_10,
	rout_sig2_10,
	iout_sig2_9,
	rout_sig2_9,
	iout_sig2_8,
	rout_sig2_8,
	b,
	a,
	iout_sig2_7,
	rout_sig2_7,
	iout_sig2_6,
	rout_sig2_6,
	iout_sig2_5,
	rout_sig2_5,
	iout_sig2_4,
	rout_sig2_4,
	iout_sig2_3,
	rout_sig2_3,
	iout_sig2_2,
	rout_sig2_2,
	iout_sig2_1,
	rout_sig2_1,
	iout_sig2_0,
	rout_sig2_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[7:0] c;
input 	[7:0] d;
input 	global_clock_enable;
output 	iout_sig2_11;
output 	iout_sig2_15;
output 	rout_sig2_11;
output 	rout_sig2_15;
output 	iout_sig2_12;
output 	rout_sig2_12;
output 	iout_sig2_13;
output 	rout_sig2_13;
output 	iout_sig2_14;
output 	rout_sig2_14;
output 	iout_sig2_10;
output 	rout_sig2_10;
output 	iout_sig2_9;
output 	rout_sig2_9;
output 	iout_sig2_8;
output 	rout_sig2_8;
input 	[7:0] b;
input 	[7:0] a;
output 	iout_sig2_7;
output 	rout_sig2_7;
output 	iout_sig2_6;
output 	rout_sig2_6;
output 	iout_sig2_5;
output 	rout_sig2_5;
output 	iout_sig2_4;
output 	rout_sig2_4;
output 	iout_sig2_3;
output 	rout_sig2_3;
output 	iout_sig2_2;
output 	rout_sig2_2;
output 	iout_sig2_1;
output 	rout_sig2_1;
output 	iout_sig2_0;
output 	rout_sig2_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~24 ;
wire \Add1~25 ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~28 ;
wire \Add1~29 ;
wire \Add1~30 ;
wire \Add1~31 ;
wire \Add1~32 ;
wire \Add1~33 ;
wire \Add1~34 ;
wire \Add1~35 ;
wire \Add1~36 ;
wire \Add1~37 ;
wire \Add1~38 ;
wire \Add1~39 ;
wire \Add1~40 ;
wire \Add1~41 ;
wire \Add1~42 ;
wire \Add1~43 ;
wire \Add1~44 ;
wire \Add1~45 ;
wire \Add1~46 ;
wire \Add1~47 ;
wire \Add1~48 ;
wire \Add1~49 ;
wire \Add1~50 ;
wire \Add1~51 ;
wire \Add1~52 ;
wire \Add1~53 ;
wire \Add1~54 ;
wire \Add1~55 ;
wire \Add1~56 ;
wire \Add1~57 ;
wire \Add1~58 ;
wire \Add1~59 ;
wire \Add1~60 ;
wire \Add1~61 ;
wire \Add1~62 ;
wire \Add1~63 ;
wire \Add1~64 ;
wire \Add1~65 ;
wire \Add1~66 ;
wire \Add1~67 ;
wire \Add1~68 ;
wire \Add1~69 ;
wire \Add1~70 ;
wire \Add1~71 ;
wire \Add0~24 ;
wire \Add0~25 ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~28 ;
wire \Add0~29 ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~32 ;
wire \Add0~33 ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~36 ;
wire \Add0~37 ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~40 ;
wire \Add0~41 ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~44 ;
wire \Add0~45 ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~48 ;
wire \Add0~49 ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~52 ;
wire \Add0~53 ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~56 ;
wire \Add0~57 ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~60 ;
wire \Add0~61 ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~64 ;
wire \Add0~65 ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~68 ;
wire \Add0~69 ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \c_reg[0]~q ;
wire \c_reg[1]~q ;
wire \c_reg[2]~q ;
wire \c_reg[3]~q ;
wire \c_reg[4]~q ;
wire \c_reg[5]~q ;
wire \c_reg[6]~q ;
wire \c_reg[7]~q ;
wire \b_reg[0]~q ;
wire \b_reg[1]~q ;
wire \b_reg[2]~q ;
wire \b_reg[3]~q ;
wire \b_reg[4]~q ;
wire \b_reg[5]~q ;
wire \b_reg[6]~q ;
wire \b_reg[7]~q ;
wire \d_reg[0]~q ;
wire \d_reg[1]~q ;
wire \d_reg[2]~q ;
wire \d_reg[3]~q ;
wire \d_reg[4]~q ;
wire \d_reg[5]~q ;
wire \d_reg[6]~q ;
wire \d_reg[7]~q ;
wire \a_reg[0]~q ;
wire \a_reg[1]~q ;
wire \a_reg[2]~q ;
wire \a_reg[3]~q ;
wire \a_reg[4]~q ;
wire \a_reg[5]~q ;
wire \a_reg[6]~q ;
wire \a_reg[7]~q ;
wire \Add1~19 ;
wire \iout_sig[11]~q ;
wire \Add1~23 ;
wire \iout_sig[15]~q ;
wire \Add0~19 ;
wire \rout_sig[11]~q ;
wire \Add0~23 ;
wire \rout_sig[15]~q ;
wire \Add1~20 ;
wire \iout_sig[12]~q ;
wire \Add0~20 ;
wire \rout_sig[12]~q ;
wire \Add1~21 ;
wire \iout_sig[13]~q ;
wire \Add0~21 ;
wire \rout_sig[13]~q ;
wire \Add1~22 ;
wire \iout_sig[14]~q ;
wire \Add0~22 ;
wire \rout_sig[14]~q ;
wire \Add1~18 ;
wire \iout_sig[10]~q ;
wire \Add0~18 ;
wire \rout_sig[10]~q ;
wire \Add1~17 ;
wire \iout_sig[9]~q ;
wire \Add0~17 ;
wire \rout_sig[9]~q ;
wire \Add1~16 ;
wire \iout_sig[8]~q ;
wire \Add0~16 ;
wire \rout_sig[8]~q ;
wire \Add1~15 ;
wire \iout_sig[7]~q ;
wire \Add0~15 ;
wire \rout_sig[7]~q ;
wire \Add1~14 ;
wire \iout_sig[6]~q ;
wire \Add0~14 ;
wire \rout_sig[6]~q ;
wire \Add1~13 ;
wire \iout_sig[5]~q ;
wire \Add0~13 ;
wire \rout_sig[5]~q ;
wire \Add1~12 ;
wire \iout_sig[4]~q ;
wire \Add0~12 ;
wire \rout_sig[4]~q ;
wire \Add1~11 ;
wire \iout_sig[3]~q ;
wire \Add0~11 ;
wire \rout_sig[3]~q ;
wire \Add1~10 ;
wire \iout_sig[2]~q ;
wire \Add0~10 ;
wire \rout_sig[2]~q ;
wire \Add1~9 ;
wire \iout_sig[1]~q ;
wire \Add0~9 ;
wire \rout_sig[1]~q ;
wire \Add1~8_resulta ;
wire \iout_sig[0]~q ;
wire \Add0~8_resulta ;
wire \rout_sig[0]~q ;

wire [63:0] \Add1~8_RESULTA_bus ;
wire [63:0] \Add0~8_RESULTA_bus ;

assign \Add1~8_resulta  = \Add1~8_RESULTA_bus [0];
assign \Add1~9  = \Add1~8_RESULTA_bus [1];
assign \Add1~10  = \Add1~8_RESULTA_bus [2];
assign \Add1~11  = \Add1~8_RESULTA_bus [3];
assign \Add1~12  = \Add1~8_RESULTA_bus [4];
assign \Add1~13  = \Add1~8_RESULTA_bus [5];
assign \Add1~14  = \Add1~8_RESULTA_bus [6];
assign \Add1~15  = \Add1~8_RESULTA_bus [7];
assign \Add1~16  = \Add1~8_RESULTA_bus [8];
assign \Add1~17  = \Add1~8_RESULTA_bus [9];
assign \Add1~18  = \Add1~8_RESULTA_bus [10];
assign \Add1~19  = \Add1~8_RESULTA_bus [11];
assign \Add1~20  = \Add1~8_RESULTA_bus [12];
assign \Add1~21  = \Add1~8_RESULTA_bus [13];
assign \Add1~22  = \Add1~8_RESULTA_bus [14];
assign \Add1~23  = \Add1~8_RESULTA_bus [15];
assign \Add1~24  = \Add1~8_RESULTA_bus [16];
assign \Add1~25  = \Add1~8_RESULTA_bus [17];
assign \Add1~26  = \Add1~8_RESULTA_bus [18];
assign \Add1~27  = \Add1~8_RESULTA_bus [19];
assign \Add1~28  = \Add1~8_RESULTA_bus [20];
assign \Add1~29  = \Add1~8_RESULTA_bus [21];
assign \Add1~30  = \Add1~8_RESULTA_bus [22];
assign \Add1~31  = \Add1~8_RESULTA_bus [23];
assign \Add1~32  = \Add1~8_RESULTA_bus [24];
assign \Add1~33  = \Add1~8_RESULTA_bus [25];
assign \Add1~34  = \Add1~8_RESULTA_bus [26];
assign \Add1~35  = \Add1~8_RESULTA_bus [27];
assign \Add1~36  = \Add1~8_RESULTA_bus [28];
assign \Add1~37  = \Add1~8_RESULTA_bus [29];
assign \Add1~38  = \Add1~8_RESULTA_bus [30];
assign \Add1~39  = \Add1~8_RESULTA_bus [31];
assign \Add1~40  = \Add1~8_RESULTA_bus [32];
assign \Add1~41  = \Add1~8_RESULTA_bus [33];
assign \Add1~42  = \Add1~8_RESULTA_bus [34];
assign \Add1~43  = \Add1~8_RESULTA_bus [35];
assign \Add1~44  = \Add1~8_RESULTA_bus [36];
assign \Add1~45  = \Add1~8_RESULTA_bus [37];
assign \Add1~46  = \Add1~8_RESULTA_bus [38];
assign \Add1~47  = \Add1~8_RESULTA_bus [39];
assign \Add1~48  = \Add1~8_RESULTA_bus [40];
assign \Add1~49  = \Add1~8_RESULTA_bus [41];
assign \Add1~50  = \Add1~8_RESULTA_bus [42];
assign \Add1~51  = \Add1~8_RESULTA_bus [43];
assign \Add1~52  = \Add1~8_RESULTA_bus [44];
assign \Add1~53  = \Add1~8_RESULTA_bus [45];
assign \Add1~54  = \Add1~8_RESULTA_bus [46];
assign \Add1~55  = \Add1~8_RESULTA_bus [47];
assign \Add1~56  = \Add1~8_RESULTA_bus [48];
assign \Add1~57  = \Add1~8_RESULTA_bus [49];
assign \Add1~58  = \Add1~8_RESULTA_bus [50];
assign \Add1~59  = \Add1~8_RESULTA_bus [51];
assign \Add1~60  = \Add1~8_RESULTA_bus [52];
assign \Add1~61  = \Add1~8_RESULTA_bus [53];
assign \Add1~62  = \Add1~8_RESULTA_bus [54];
assign \Add1~63  = \Add1~8_RESULTA_bus [55];
assign \Add1~64  = \Add1~8_RESULTA_bus [56];
assign \Add1~65  = \Add1~8_RESULTA_bus [57];
assign \Add1~66  = \Add1~8_RESULTA_bus [58];
assign \Add1~67  = \Add1~8_RESULTA_bus [59];
assign \Add1~68  = \Add1~8_RESULTA_bus [60];
assign \Add1~69  = \Add1~8_RESULTA_bus [61];
assign \Add1~70  = \Add1~8_RESULTA_bus [62];
assign \Add1~71  = \Add1~8_RESULTA_bus [63];

assign \Add0~8_resulta  = \Add0~8_RESULTA_bus [0];
assign \Add0~9  = \Add0~8_RESULTA_bus [1];
assign \Add0~10  = \Add0~8_RESULTA_bus [2];
assign \Add0~11  = \Add0~8_RESULTA_bus [3];
assign \Add0~12  = \Add0~8_RESULTA_bus [4];
assign \Add0~13  = \Add0~8_RESULTA_bus [5];
assign \Add0~14  = \Add0~8_RESULTA_bus [6];
assign \Add0~15  = \Add0~8_RESULTA_bus [7];
assign \Add0~16  = \Add0~8_RESULTA_bus [8];
assign \Add0~17  = \Add0~8_RESULTA_bus [9];
assign \Add0~18  = \Add0~8_RESULTA_bus [10];
assign \Add0~19  = \Add0~8_RESULTA_bus [11];
assign \Add0~20  = \Add0~8_RESULTA_bus [12];
assign \Add0~21  = \Add0~8_RESULTA_bus [13];
assign \Add0~22  = \Add0~8_RESULTA_bus [14];
assign \Add0~23  = \Add0~8_RESULTA_bus [15];
assign \Add0~24  = \Add0~8_RESULTA_bus [16];
assign \Add0~25  = \Add0~8_RESULTA_bus [17];
assign \Add0~26  = \Add0~8_RESULTA_bus [18];
assign \Add0~27  = \Add0~8_RESULTA_bus [19];
assign \Add0~28  = \Add0~8_RESULTA_bus [20];
assign \Add0~29  = \Add0~8_RESULTA_bus [21];
assign \Add0~30  = \Add0~8_RESULTA_bus [22];
assign \Add0~31  = \Add0~8_RESULTA_bus [23];
assign \Add0~32  = \Add0~8_RESULTA_bus [24];
assign \Add0~33  = \Add0~8_RESULTA_bus [25];
assign \Add0~34  = \Add0~8_RESULTA_bus [26];
assign \Add0~35  = \Add0~8_RESULTA_bus [27];
assign \Add0~36  = \Add0~8_RESULTA_bus [28];
assign \Add0~37  = \Add0~8_RESULTA_bus [29];
assign \Add0~38  = \Add0~8_RESULTA_bus [30];
assign \Add0~39  = \Add0~8_RESULTA_bus [31];
assign \Add0~40  = \Add0~8_RESULTA_bus [32];
assign \Add0~41  = \Add0~8_RESULTA_bus [33];
assign \Add0~42  = \Add0~8_RESULTA_bus [34];
assign \Add0~43  = \Add0~8_RESULTA_bus [35];
assign \Add0~44  = \Add0~8_RESULTA_bus [36];
assign \Add0~45  = \Add0~8_RESULTA_bus [37];
assign \Add0~46  = \Add0~8_RESULTA_bus [38];
assign \Add0~47  = \Add0~8_RESULTA_bus [39];
assign \Add0~48  = \Add0~8_RESULTA_bus [40];
assign \Add0~49  = \Add0~8_RESULTA_bus [41];
assign \Add0~50  = \Add0~8_RESULTA_bus [42];
assign \Add0~51  = \Add0~8_RESULTA_bus [43];
assign \Add0~52  = \Add0~8_RESULTA_bus [44];
assign \Add0~53  = \Add0~8_RESULTA_bus [45];
assign \Add0~54  = \Add0~8_RESULTA_bus [46];
assign \Add0~55  = \Add0~8_RESULTA_bus [47];
assign \Add0~56  = \Add0~8_RESULTA_bus [48];
assign \Add0~57  = \Add0~8_RESULTA_bus [49];
assign \Add0~58  = \Add0~8_RESULTA_bus [50];
assign \Add0~59  = \Add0~8_RESULTA_bus [51];
assign \Add0~60  = \Add0~8_RESULTA_bus [52];
assign \Add0~61  = \Add0~8_RESULTA_bus [53];
assign \Add0~62  = \Add0~8_RESULTA_bus [54];
assign \Add0~63  = \Add0~8_RESULTA_bus [55];
assign \Add0~64  = \Add0~8_RESULTA_bus [56];
assign \Add0~65  = \Add0~8_RESULTA_bus [57];
assign \Add0~66  = \Add0~8_RESULTA_bus [58];
assign \Add0~67  = \Add0~8_RESULTA_bus [59];
assign \Add0~68  = \Add0~8_RESULTA_bus [60];
assign \Add0~69  = \Add0~8_RESULTA_bus [61];
assign \Add0~70  = \Add0~8_RESULTA_bus [62];
assign \Add0~71  = \Add0~8_RESULTA_bus [63];

dffeas \iout_sig2[11] (
	.clk(clk),
	.d(\iout_sig[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_11),
	.prn(vcc));
defparam \iout_sig2[11] .is_wysiwyg = "true";
defparam \iout_sig2[11] .power_up = "low";

dffeas \iout_sig2[15] (
	.clk(clk),
	.d(\iout_sig[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_15),
	.prn(vcc));
defparam \iout_sig2[15] .is_wysiwyg = "true";
defparam \iout_sig2[15] .power_up = "low";

dffeas \rout_sig2[11] (
	.clk(clk),
	.d(\rout_sig[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_11),
	.prn(vcc));
defparam \rout_sig2[11] .is_wysiwyg = "true";
defparam \rout_sig2[11] .power_up = "low";

dffeas \rout_sig2[15] (
	.clk(clk),
	.d(\rout_sig[15]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_15),
	.prn(vcc));
defparam \rout_sig2[15] .is_wysiwyg = "true";
defparam \rout_sig2[15] .power_up = "low";

dffeas \iout_sig2[12] (
	.clk(clk),
	.d(\iout_sig[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_12),
	.prn(vcc));
defparam \iout_sig2[12] .is_wysiwyg = "true";
defparam \iout_sig2[12] .power_up = "low";

dffeas \rout_sig2[12] (
	.clk(clk),
	.d(\rout_sig[12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_12),
	.prn(vcc));
defparam \rout_sig2[12] .is_wysiwyg = "true";
defparam \rout_sig2[12] .power_up = "low";

dffeas \iout_sig2[13] (
	.clk(clk),
	.d(\iout_sig[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_13),
	.prn(vcc));
defparam \iout_sig2[13] .is_wysiwyg = "true";
defparam \iout_sig2[13] .power_up = "low";

dffeas \rout_sig2[13] (
	.clk(clk),
	.d(\rout_sig[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_13),
	.prn(vcc));
defparam \rout_sig2[13] .is_wysiwyg = "true";
defparam \rout_sig2[13] .power_up = "low";

dffeas \iout_sig2[14] (
	.clk(clk),
	.d(\iout_sig[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_14),
	.prn(vcc));
defparam \iout_sig2[14] .is_wysiwyg = "true";
defparam \iout_sig2[14] .power_up = "low";

dffeas \rout_sig2[14] (
	.clk(clk),
	.d(\rout_sig[14]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_14),
	.prn(vcc));
defparam \rout_sig2[14] .is_wysiwyg = "true";
defparam \rout_sig2[14] .power_up = "low";

dffeas \iout_sig2[10] (
	.clk(clk),
	.d(\iout_sig[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_10),
	.prn(vcc));
defparam \iout_sig2[10] .is_wysiwyg = "true";
defparam \iout_sig2[10] .power_up = "low";

dffeas \rout_sig2[10] (
	.clk(clk),
	.d(\rout_sig[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_10),
	.prn(vcc));
defparam \rout_sig2[10] .is_wysiwyg = "true";
defparam \rout_sig2[10] .power_up = "low";

dffeas \iout_sig2[9] (
	.clk(clk),
	.d(\iout_sig[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_9),
	.prn(vcc));
defparam \iout_sig2[9] .is_wysiwyg = "true";
defparam \iout_sig2[9] .power_up = "low";

dffeas \rout_sig2[9] (
	.clk(clk),
	.d(\rout_sig[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_9),
	.prn(vcc));
defparam \rout_sig2[9] .is_wysiwyg = "true";
defparam \rout_sig2[9] .power_up = "low";

dffeas \iout_sig2[8] (
	.clk(clk),
	.d(\iout_sig[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_8),
	.prn(vcc));
defparam \iout_sig2[8] .is_wysiwyg = "true";
defparam \iout_sig2[8] .power_up = "low";

dffeas \rout_sig2[8] (
	.clk(clk),
	.d(\rout_sig[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_8),
	.prn(vcc));
defparam \rout_sig2[8] .is_wysiwyg = "true";
defparam \rout_sig2[8] .power_up = "low";

dffeas \iout_sig2[7] (
	.clk(clk),
	.d(\iout_sig[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_7),
	.prn(vcc));
defparam \iout_sig2[7] .is_wysiwyg = "true";
defparam \iout_sig2[7] .power_up = "low";

dffeas \rout_sig2[7] (
	.clk(clk),
	.d(\rout_sig[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_7),
	.prn(vcc));
defparam \rout_sig2[7] .is_wysiwyg = "true";
defparam \rout_sig2[7] .power_up = "low";

dffeas \iout_sig2[6] (
	.clk(clk),
	.d(\iout_sig[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_6),
	.prn(vcc));
defparam \iout_sig2[6] .is_wysiwyg = "true";
defparam \iout_sig2[6] .power_up = "low";

dffeas \rout_sig2[6] (
	.clk(clk),
	.d(\rout_sig[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_6),
	.prn(vcc));
defparam \rout_sig2[6] .is_wysiwyg = "true";
defparam \rout_sig2[6] .power_up = "low";

dffeas \iout_sig2[5] (
	.clk(clk),
	.d(\iout_sig[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_5),
	.prn(vcc));
defparam \iout_sig2[5] .is_wysiwyg = "true";
defparam \iout_sig2[5] .power_up = "low";

dffeas \rout_sig2[5] (
	.clk(clk),
	.d(\rout_sig[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_5),
	.prn(vcc));
defparam \rout_sig2[5] .is_wysiwyg = "true";
defparam \rout_sig2[5] .power_up = "low";

dffeas \iout_sig2[4] (
	.clk(clk),
	.d(\iout_sig[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_4),
	.prn(vcc));
defparam \iout_sig2[4] .is_wysiwyg = "true";
defparam \iout_sig2[4] .power_up = "low";

dffeas \rout_sig2[4] (
	.clk(clk),
	.d(\rout_sig[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_4),
	.prn(vcc));
defparam \rout_sig2[4] .is_wysiwyg = "true";
defparam \rout_sig2[4] .power_up = "low";

dffeas \iout_sig2[3] (
	.clk(clk),
	.d(\iout_sig[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_3),
	.prn(vcc));
defparam \iout_sig2[3] .is_wysiwyg = "true";
defparam \iout_sig2[3] .power_up = "low";

dffeas \rout_sig2[3] (
	.clk(clk),
	.d(\rout_sig[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_3),
	.prn(vcc));
defparam \rout_sig2[3] .is_wysiwyg = "true";
defparam \rout_sig2[3] .power_up = "low";

dffeas \iout_sig2[2] (
	.clk(clk),
	.d(\iout_sig[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_2),
	.prn(vcc));
defparam \iout_sig2[2] .is_wysiwyg = "true";
defparam \iout_sig2[2] .power_up = "low";

dffeas \rout_sig2[2] (
	.clk(clk),
	.d(\rout_sig[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_2),
	.prn(vcc));
defparam \rout_sig2[2] .is_wysiwyg = "true";
defparam \rout_sig2[2] .power_up = "low";

dffeas \iout_sig2[1] (
	.clk(clk),
	.d(\iout_sig[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_1),
	.prn(vcc));
defparam \iout_sig2[1] .is_wysiwyg = "true";
defparam \iout_sig2[1] .power_up = "low";

dffeas \rout_sig2[1] (
	.clk(clk),
	.d(\rout_sig[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_1),
	.prn(vcc));
defparam \rout_sig2[1] .is_wysiwyg = "true";
defparam \rout_sig2[1] .power_up = "low";

dffeas \iout_sig2[0] (
	.clk(clk),
	.d(\iout_sig[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(iout_sig2_0),
	.prn(vcc));
defparam \iout_sig2[0] .is_wysiwyg = "true";
defparam \iout_sig2[0] .power_up = "low";

dffeas \rout_sig2[0] (
	.clk(clk),
	.d(\rout_sig[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rout_sig2_0),
	.prn(vcc));
defparam \rout_sig2[0] .is_wysiwyg = "true";
defparam \rout_sig2[0] .power_up = "low";

dffeas \c_reg[0] (
	.clk(clk),
	.d(c[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[0]~q ),
	.prn(vcc));
defparam \c_reg[0] .is_wysiwyg = "true";
defparam \c_reg[0] .power_up = "low";

dffeas \c_reg[1] (
	.clk(clk),
	.d(c[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[1]~q ),
	.prn(vcc));
defparam \c_reg[1] .is_wysiwyg = "true";
defparam \c_reg[1] .power_up = "low";

dffeas \c_reg[2] (
	.clk(clk),
	.d(c[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[2]~q ),
	.prn(vcc));
defparam \c_reg[2] .is_wysiwyg = "true";
defparam \c_reg[2] .power_up = "low";

dffeas \c_reg[3] (
	.clk(clk),
	.d(c[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[3]~q ),
	.prn(vcc));
defparam \c_reg[3] .is_wysiwyg = "true";
defparam \c_reg[3] .power_up = "low";

dffeas \c_reg[4] (
	.clk(clk),
	.d(c[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[4]~q ),
	.prn(vcc));
defparam \c_reg[4] .is_wysiwyg = "true";
defparam \c_reg[4] .power_up = "low";

dffeas \c_reg[5] (
	.clk(clk),
	.d(c[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[5]~q ),
	.prn(vcc));
defparam \c_reg[5] .is_wysiwyg = "true";
defparam \c_reg[5] .power_up = "low";

dffeas \c_reg[6] (
	.clk(clk),
	.d(c[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[6]~q ),
	.prn(vcc));
defparam \c_reg[6] .is_wysiwyg = "true";
defparam \c_reg[6] .power_up = "low";

dffeas \c_reg[7] (
	.clk(clk),
	.d(c[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\c_reg[7]~q ),
	.prn(vcc));
defparam \c_reg[7] .is_wysiwyg = "true";
defparam \c_reg[7] .power_up = "low";

dffeas \b_reg[0] (
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[0]~q ),
	.prn(vcc));
defparam \b_reg[0] .is_wysiwyg = "true";
defparam \b_reg[0] .power_up = "low";

dffeas \b_reg[1] (
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[1]~q ),
	.prn(vcc));
defparam \b_reg[1] .is_wysiwyg = "true";
defparam \b_reg[1] .power_up = "low";

dffeas \b_reg[2] (
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[2]~q ),
	.prn(vcc));
defparam \b_reg[2] .is_wysiwyg = "true";
defparam \b_reg[2] .power_up = "low";

dffeas \b_reg[3] (
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[3]~q ),
	.prn(vcc));
defparam \b_reg[3] .is_wysiwyg = "true";
defparam \b_reg[3] .power_up = "low";

dffeas \b_reg[4] (
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[4]~q ),
	.prn(vcc));
defparam \b_reg[4] .is_wysiwyg = "true";
defparam \b_reg[4] .power_up = "low";

dffeas \b_reg[5] (
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[5]~q ),
	.prn(vcc));
defparam \b_reg[5] .is_wysiwyg = "true";
defparam \b_reg[5] .power_up = "low";

dffeas \b_reg[6] (
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[6]~q ),
	.prn(vcc));
defparam \b_reg[6] .is_wysiwyg = "true";
defparam \b_reg[6] .power_up = "low";

dffeas \b_reg[7] (
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\b_reg[7]~q ),
	.prn(vcc));
defparam \b_reg[7] .is_wysiwyg = "true";
defparam \b_reg[7] .power_up = "low";

dffeas \d_reg[0] (
	.clk(clk),
	.d(d[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[0]~q ),
	.prn(vcc));
defparam \d_reg[0] .is_wysiwyg = "true";
defparam \d_reg[0] .power_up = "low";

dffeas \d_reg[1] (
	.clk(clk),
	.d(d[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[1]~q ),
	.prn(vcc));
defparam \d_reg[1] .is_wysiwyg = "true";
defparam \d_reg[1] .power_up = "low";

dffeas \d_reg[2] (
	.clk(clk),
	.d(d[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[2]~q ),
	.prn(vcc));
defparam \d_reg[2] .is_wysiwyg = "true";
defparam \d_reg[2] .power_up = "low";

dffeas \d_reg[3] (
	.clk(clk),
	.d(d[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[3]~q ),
	.prn(vcc));
defparam \d_reg[3] .is_wysiwyg = "true";
defparam \d_reg[3] .power_up = "low";

dffeas \d_reg[4] (
	.clk(clk),
	.d(d[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[4]~q ),
	.prn(vcc));
defparam \d_reg[4] .is_wysiwyg = "true";
defparam \d_reg[4] .power_up = "low";

dffeas \d_reg[5] (
	.clk(clk),
	.d(d[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[5]~q ),
	.prn(vcc));
defparam \d_reg[5] .is_wysiwyg = "true";
defparam \d_reg[5] .power_up = "low";

dffeas \d_reg[6] (
	.clk(clk),
	.d(d[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[6]~q ),
	.prn(vcc));
defparam \d_reg[6] .is_wysiwyg = "true";
defparam \d_reg[6] .power_up = "low";

dffeas \d_reg[7] (
	.clk(clk),
	.d(d[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\d_reg[7]~q ),
	.prn(vcc));
defparam \d_reg[7] .is_wysiwyg = "true";
defparam \d_reg[7] .power_up = "low";

dffeas \a_reg[0] (
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[0]~q ),
	.prn(vcc));
defparam \a_reg[0] .is_wysiwyg = "true";
defparam \a_reg[0] .power_up = "low";

dffeas \a_reg[1] (
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[1]~q ),
	.prn(vcc));
defparam \a_reg[1] .is_wysiwyg = "true";
defparam \a_reg[1] .power_up = "low";

dffeas \a_reg[2] (
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[2]~q ),
	.prn(vcc));
defparam \a_reg[2] .is_wysiwyg = "true";
defparam \a_reg[2] .power_up = "low";

dffeas \a_reg[3] (
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[3]~q ),
	.prn(vcc));
defparam \a_reg[3] .is_wysiwyg = "true";
defparam \a_reg[3] .power_up = "low";

dffeas \a_reg[4] (
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[4]~q ),
	.prn(vcc));
defparam \a_reg[4] .is_wysiwyg = "true";
defparam \a_reg[4] .power_up = "low";

dffeas \a_reg[5] (
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[5]~q ),
	.prn(vcc));
defparam \a_reg[5] .is_wysiwyg = "true";
defparam \a_reg[5] .power_up = "low";

dffeas \a_reg[6] (
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[6]~q ),
	.prn(vcc));
defparam \a_reg[6] .is_wysiwyg = "true";
defparam \a_reg[6] .power_up = "low";

dffeas \a_reg[7] (
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\a_reg[7]~q ),
	.prn(vcc));
defparam \a_reg[7] .is_wysiwyg = "true";
defparam \a_reg[7] .power_up = "low";

cyclonev_mac \Add1~8 (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\c_reg[7]~q ,\c_reg[6]~q ,\c_reg[5]~q ,\c_reg[4]~q ,\c_reg[3]~q ,\c_reg[2]~q ,\c_reg[1]~q ,\c_reg[0]~q }),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\b_reg[7]~q ,\b_reg[6]~q ,\b_reg[5]~q ,\b_reg[4]~q ,\b_reg[3]~q ,\b_reg[2]~q ,\b_reg[1]~q ,\b_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_reg[7]~q ,\d_reg[6]~q ,\d_reg[5]~q ,\d_reg[4]~q ,\d_reg[3]~q ,\d_reg[2]~q ,\d_reg[1]~q ,\d_reg[0]~q }),
	.by({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\a_reg[7]~q ,\a_reg[6]~q ,\a_reg[5]~q ,\a_reg[4]~q ,\a_reg[3]~q ,\a_reg[2]~q ,\a_reg[1]~q ,\a_reg[0]~q }),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Add1~8_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Add1~8 .accumulate_clock = "none";
defparam \Add1~8 .ax_clock = "none";
defparam \Add1~8 .ax_width = 8;
defparam \Add1~8 .ay_scan_in_clock = "none";
defparam \Add1~8 .ay_scan_in_width = 8;
defparam \Add1~8 .ay_use_scan_in = "false";
defparam \Add1~8 .az_clock = "none";
defparam \Add1~8 .bx_clock = "none";
defparam \Add1~8 .bx_width = 8;
defparam \Add1~8 .by_clock = "none";
defparam \Add1~8 .by_use_scan_in = "false";
defparam \Add1~8 .by_width = 8;
defparam \Add1~8 .bz_clock = "none";
defparam \Add1~8 .coef_a_0 = 0;
defparam \Add1~8 .coef_a_1 = 0;
defparam \Add1~8 .coef_a_2 = 0;
defparam \Add1~8 .coef_a_3 = 0;
defparam \Add1~8 .coef_a_4 = 0;
defparam \Add1~8 .coef_a_5 = 0;
defparam \Add1~8 .coef_a_6 = 0;
defparam \Add1~8 .coef_a_7 = 0;
defparam \Add1~8 .coef_b_0 = 0;
defparam \Add1~8 .coef_b_1 = 0;
defparam \Add1~8 .coef_b_2 = 0;
defparam \Add1~8 .coef_b_3 = 0;
defparam \Add1~8 .coef_b_4 = 0;
defparam \Add1~8 .coef_b_5 = 0;
defparam \Add1~8 .coef_b_6 = 0;
defparam \Add1~8 .coef_b_7 = 0;
defparam \Add1~8 .coef_sel_a_clock = "none";
defparam \Add1~8 .coef_sel_b_clock = "none";
defparam \Add1~8 .delay_scan_out_ay = "false";
defparam \Add1~8 .delay_scan_out_by = "false";
defparam \Add1~8 .enable_double_accum = "false";
defparam \Add1~8 .load_const_clock = "none";
defparam \Add1~8 .load_const_value = 0;
defparam \Add1~8 .mode_sub_location = 0;
defparam \Add1~8 .negate_clock = "none";
defparam \Add1~8 .operand_source_max = "input";
defparam \Add1~8 .operand_source_may = "input";
defparam \Add1~8 .operand_source_mbx = "input";
defparam \Add1~8 .operand_source_mby = "input";
defparam \Add1~8 .operation_mode = "m18x18_sumof2";
defparam \Add1~8 .output_clock = "none";
defparam \Add1~8 .preadder_subtract_a = "false";
defparam \Add1~8 .preadder_subtract_b = "false";
defparam \Add1~8 .result_a_width = 64;
defparam \Add1~8 .signed_max = "true";
defparam \Add1~8 .signed_may = "true";
defparam \Add1~8 .signed_mbx = "true";
defparam \Add1~8 .signed_mby = "true";
defparam \Add1~8 .sub_clock = "none";
defparam \Add1~8 .use_chainadder = "false";

dffeas \iout_sig[11] (
	.clk(clk),
	.d(\Add1~19 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[11]~q ),
	.prn(vcc));
defparam \iout_sig[11] .is_wysiwyg = "true";
defparam \iout_sig[11] .power_up = "low";

dffeas \iout_sig[15] (
	.clk(clk),
	.d(\Add1~23 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[15]~q ),
	.prn(vcc));
defparam \iout_sig[15] .is_wysiwyg = "true";
defparam \iout_sig[15] .power_up = "low";

cyclonev_mac \Add0~8 (
	.sub(vcc),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\d_reg[7]~q ,\d_reg[6]~q ,\d_reg[5]~q ,\d_reg[4]~q ,\d_reg[3]~q ,\d_reg[2]~q ,\d_reg[1]~q ,\d_reg[0]~q }),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\b_reg[7]~q ,\b_reg[6]~q ,\b_reg[5]~q ,\b_reg[4]~q ,\b_reg[3]~q ,\b_reg[2]~q ,\b_reg[1]~q ,\b_reg[0]~q }),
	.az(26'b00000000000000000000000000),
	.bx({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\c_reg[7]~q ,\c_reg[6]~q ,\c_reg[5]~q ,\c_reg[4]~q ,\c_reg[3]~q ,\c_reg[2]~q ,\c_reg[1]~q ,\c_reg[0]~q }),
	.by({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\a_reg[7]~q ,\a_reg[6]~q ,\a_reg[5]~q ,\a_reg[4]~q ,\a_reg[3]~q ,\a_reg[2]~q ,\a_reg[1]~q ,\a_reg[0]~q }),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Add0~8_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Add0~8 .accumulate_clock = "none";
defparam \Add0~8 .ax_clock = "none";
defparam \Add0~8 .ax_width = 8;
defparam \Add0~8 .ay_scan_in_clock = "none";
defparam \Add0~8 .ay_scan_in_width = 8;
defparam \Add0~8 .ay_use_scan_in = "false";
defparam \Add0~8 .az_clock = "none";
defparam \Add0~8 .bx_clock = "none";
defparam \Add0~8 .bx_width = 8;
defparam \Add0~8 .by_clock = "none";
defparam \Add0~8 .by_use_scan_in = "false";
defparam \Add0~8 .by_width = 8;
defparam \Add0~8 .bz_clock = "none";
defparam \Add0~8 .coef_a_0 = 0;
defparam \Add0~8 .coef_a_1 = 0;
defparam \Add0~8 .coef_a_2 = 0;
defparam \Add0~8 .coef_a_3 = 0;
defparam \Add0~8 .coef_a_4 = 0;
defparam \Add0~8 .coef_a_5 = 0;
defparam \Add0~8 .coef_a_6 = 0;
defparam \Add0~8 .coef_a_7 = 0;
defparam \Add0~8 .coef_b_0 = 0;
defparam \Add0~8 .coef_b_1 = 0;
defparam \Add0~8 .coef_b_2 = 0;
defparam \Add0~8 .coef_b_3 = 0;
defparam \Add0~8 .coef_b_4 = 0;
defparam \Add0~8 .coef_b_5 = 0;
defparam \Add0~8 .coef_b_6 = 0;
defparam \Add0~8 .coef_b_7 = 0;
defparam \Add0~8 .coef_sel_a_clock = "none";
defparam \Add0~8 .coef_sel_b_clock = "none";
defparam \Add0~8 .delay_scan_out_ay = "false";
defparam \Add0~8 .delay_scan_out_by = "false";
defparam \Add0~8 .enable_double_accum = "false";
defparam \Add0~8 .load_const_clock = "none";
defparam \Add0~8 .load_const_value = 0;
defparam \Add0~8 .mode_sub_location = 0;
defparam \Add0~8 .negate_clock = "none";
defparam \Add0~8 .operand_source_max = "input";
defparam \Add0~8 .operand_source_may = "input";
defparam \Add0~8 .operand_source_mbx = "input";
defparam \Add0~8 .operand_source_mby = "input";
defparam \Add0~8 .operation_mode = "m18x18_sumof2";
defparam \Add0~8 .output_clock = "none";
defparam \Add0~8 .preadder_subtract_a = "false";
defparam \Add0~8 .preadder_subtract_b = "false";
defparam \Add0~8 .result_a_width = 64;
defparam \Add0~8 .signed_max = "true";
defparam \Add0~8 .signed_may = "true";
defparam \Add0~8 .signed_mbx = "true";
defparam \Add0~8 .signed_mby = "true";
defparam \Add0~8 .sub_clock = "none";
defparam \Add0~8 .use_chainadder = "false";

dffeas \rout_sig[11] (
	.clk(clk),
	.d(\Add0~19 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[11]~q ),
	.prn(vcc));
defparam \rout_sig[11] .is_wysiwyg = "true";
defparam \rout_sig[11] .power_up = "low";

dffeas \rout_sig[15] (
	.clk(clk),
	.d(\Add0~23 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[15]~q ),
	.prn(vcc));
defparam \rout_sig[15] .is_wysiwyg = "true";
defparam \rout_sig[15] .power_up = "low";

dffeas \iout_sig[12] (
	.clk(clk),
	.d(\Add1~20 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[12]~q ),
	.prn(vcc));
defparam \iout_sig[12] .is_wysiwyg = "true";
defparam \iout_sig[12] .power_up = "low";

dffeas \rout_sig[12] (
	.clk(clk),
	.d(\Add0~20 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[12]~q ),
	.prn(vcc));
defparam \rout_sig[12] .is_wysiwyg = "true";
defparam \rout_sig[12] .power_up = "low";

dffeas \iout_sig[13] (
	.clk(clk),
	.d(\Add1~21 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[13]~q ),
	.prn(vcc));
defparam \iout_sig[13] .is_wysiwyg = "true";
defparam \iout_sig[13] .power_up = "low";

dffeas \rout_sig[13] (
	.clk(clk),
	.d(\Add0~21 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[13]~q ),
	.prn(vcc));
defparam \rout_sig[13] .is_wysiwyg = "true";
defparam \rout_sig[13] .power_up = "low";

dffeas \iout_sig[14] (
	.clk(clk),
	.d(\Add1~22 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[14]~q ),
	.prn(vcc));
defparam \iout_sig[14] .is_wysiwyg = "true";
defparam \iout_sig[14] .power_up = "low";

dffeas \rout_sig[14] (
	.clk(clk),
	.d(\Add0~22 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[14]~q ),
	.prn(vcc));
defparam \rout_sig[14] .is_wysiwyg = "true";
defparam \rout_sig[14] .power_up = "low";

dffeas \iout_sig[10] (
	.clk(clk),
	.d(\Add1~18 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[10]~q ),
	.prn(vcc));
defparam \iout_sig[10] .is_wysiwyg = "true";
defparam \iout_sig[10] .power_up = "low";

dffeas \rout_sig[10] (
	.clk(clk),
	.d(\Add0~18 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[10]~q ),
	.prn(vcc));
defparam \rout_sig[10] .is_wysiwyg = "true";
defparam \rout_sig[10] .power_up = "low";

dffeas \iout_sig[9] (
	.clk(clk),
	.d(\Add1~17 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[9]~q ),
	.prn(vcc));
defparam \iout_sig[9] .is_wysiwyg = "true";
defparam \iout_sig[9] .power_up = "low";

dffeas \rout_sig[9] (
	.clk(clk),
	.d(\Add0~17 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[9]~q ),
	.prn(vcc));
defparam \rout_sig[9] .is_wysiwyg = "true";
defparam \rout_sig[9] .power_up = "low";

dffeas \iout_sig[8] (
	.clk(clk),
	.d(\Add1~16 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[8]~q ),
	.prn(vcc));
defparam \iout_sig[8] .is_wysiwyg = "true";
defparam \iout_sig[8] .power_up = "low";

dffeas \rout_sig[8] (
	.clk(clk),
	.d(\Add0~16 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[8]~q ),
	.prn(vcc));
defparam \rout_sig[8] .is_wysiwyg = "true";
defparam \rout_sig[8] .power_up = "low";

dffeas \iout_sig[7] (
	.clk(clk),
	.d(\Add1~15 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[7]~q ),
	.prn(vcc));
defparam \iout_sig[7] .is_wysiwyg = "true";
defparam \iout_sig[7] .power_up = "low";

dffeas \rout_sig[7] (
	.clk(clk),
	.d(\Add0~15 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[7]~q ),
	.prn(vcc));
defparam \rout_sig[7] .is_wysiwyg = "true";
defparam \rout_sig[7] .power_up = "low";

dffeas \iout_sig[6] (
	.clk(clk),
	.d(\Add1~14 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[6]~q ),
	.prn(vcc));
defparam \iout_sig[6] .is_wysiwyg = "true";
defparam \iout_sig[6] .power_up = "low";

dffeas \rout_sig[6] (
	.clk(clk),
	.d(\Add0~14 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[6]~q ),
	.prn(vcc));
defparam \rout_sig[6] .is_wysiwyg = "true";
defparam \rout_sig[6] .power_up = "low";

dffeas \iout_sig[5] (
	.clk(clk),
	.d(\Add1~13 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[5]~q ),
	.prn(vcc));
defparam \iout_sig[5] .is_wysiwyg = "true";
defparam \iout_sig[5] .power_up = "low";

dffeas \rout_sig[5] (
	.clk(clk),
	.d(\Add0~13 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[5]~q ),
	.prn(vcc));
defparam \rout_sig[5] .is_wysiwyg = "true";
defparam \rout_sig[5] .power_up = "low";

dffeas \iout_sig[4] (
	.clk(clk),
	.d(\Add1~12 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[4]~q ),
	.prn(vcc));
defparam \iout_sig[4] .is_wysiwyg = "true";
defparam \iout_sig[4] .power_up = "low";

dffeas \rout_sig[4] (
	.clk(clk),
	.d(\Add0~12 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[4]~q ),
	.prn(vcc));
defparam \rout_sig[4] .is_wysiwyg = "true";
defparam \rout_sig[4] .power_up = "low";

dffeas \iout_sig[3] (
	.clk(clk),
	.d(\Add1~11 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[3]~q ),
	.prn(vcc));
defparam \iout_sig[3] .is_wysiwyg = "true";
defparam \iout_sig[3] .power_up = "low";

dffeas \rout_sig[3] (
	.clk(clk),
	.d(\Add0~11 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[3]~q ),
	.prn(vcc));
defparam \rout_sig[3] .is_wysiwyg = "true";
defparam \rout_sig[3] .power_up = "low";

dffeas \iout_sig[2] (
	.clk(clk),
	.d(\Add1~10 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[2]~q ),
	.prn(vcc));
defparam \iout_sig[2] .is_wysiwyg = "true";
defparam \iout_sig[2] .power_up = "low";

dffeas \rout_sig[2] (
	.clk(clk),
	.d(\Add0~10 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[2]~q ),
	.prn(vcc));
defparam \rout_sig[2] .is_wysiwyg = "true";
defparam \rout_sig[2] .power_up = "low";

dffeas \iout_sig[1] (
	.clk(clk),
	.d(\Add1~9 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[1]~q ),
	.prn(vcc));
defparam \iout_sig[1] .is_wysiwyg = "true";
defparam \iout_sig[1] .power_up = "low";

dffeas \rout_sig[1] (
	.clk(clk),
	.d(\Add0~9 ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[1]~q ),
	.prn(vcc));
defparam \rout_sig[1] .is_wysiwyg = "true";
defparam \rout_sig[1] .power_up = "low";

dffeas \iout_sig[0] (
	.clk(clk),
	.d(\Add1~8_resulta ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\iout_sig[0]~q ),
	.prn(vcc));
defparam \iout_sig[0] .is_wysiwyg = "true";
defparam \iout_sig[0] .power_up = "low";

dffeas \rout_sig[0] (
	.clk(clk),
	.d(\Add0~8_resulta ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\rout_sig[0]~q ),
	.prn(vcc));
defparam \rout_sig[0] .is_wysiwyg = "true";
defparam \rout_sig[0] .power_up = "low";

endmodule

module IFFT_asj_fft_pround_4 (
	global_clock_enable,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_5 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_r_tmp_8(result_r_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_r_tmp_7(result_r_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_5 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_8gj_4 auto_generated(
	.clken(clken),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_r_tmp_11(result_r_tmp_11),
	.result_r_tmp_15(result_r_tmp_15),
	.result_r_tmp_12(result_r_tmp_12),
	.result_r_tmp_13(result_r_tmp_13),
	.result_r_tmp_14(result_r_tmp_14),
	.result_r_tmp_10(result_r_tmp_10),
	.result_r_tmp_9(result_r_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_r_tmp_8(result_r_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_r_tmp_7(result_r_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_r_tmp_6(result_r_tmp_6),
	.result_r_tmp_5(result_r_tmp_5),
	.result_r_tmp_4(result_r_tmp_4),
	.result_r_tmp_3(result_r_tmp_3),
	.result_r_tmp_2(result_r_tmp_2),
	.result_r_tmp_1(result_r_tmp_1),
	.result_r_tmp_0(result_r_tmp_0),
	.clock(clock));

endmodule

module IFFT_add_sub_8gj_4 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_r_tmp_11,
	result_r_tmp_15,
	result_r_tmp_12,
	result_r_tmp_13,
	result_r_tmp_14,
	result_r_tmp_10,
	result_r_tmp_9,
	pipeline_dffe_10,
	result_r_tmp_8,
	pipeline_dffe_9,
	result_r_tmp_7,
	pipeline_dffe_8,
	result_r_tmp_6,
	result_r_tmp_5,
	result_r_tmp_4,
	result_r_tmp_3,
	result_r_tmp_2,
	result_r_tmp_1,
	result_r_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_r_tmp_11;
input 	result_r_tmp_15;
input 	result_r_tmp_12;
input 	result_r_tmp_13;
input 	result_r_tmp_14;
input 	result_r_tmp_10;
input 	result_r_tmp_9;
output 	pipeline_dffe_10;
input 	result_r_tmp_8;
output 	pipeline_dffe_9;
input 	result_r_tmp_7;
output 	pipeline_dffe_8;
input 	result_r_tmp_6;
input 	result_r_tmp_5;
input 	result_r_tmp_4;
input 	result_r_tmp_3;
input 	result_r_tmp_2;
input 	result_r_tmp_1;
input 	result_r_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_r_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_5 (
	global_clock_enable,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_6 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_i_tmp_8(result_i_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_i_tmp_7(result_i_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_6 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_8gj_5 auto_generated(
	.clken(clken),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.result_i_tmp_11(result_i_tmp_11),
	.result_i_tmp_15(result_i_tmp_15),
	.result_i_tmp_12(result_i_tmp_12),
	.result_i_tmp_13(result_i_tmp_13),
	.result_i_tmp_14(result_i_tmp_14),
	.result_i_tmp_10(result_i_tmp_10),
	.result_i_tmp_9(result_i_tmp_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.result_i_tmp_8(result_i_tmp_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.result_i_tmp_7(result_i_tmp_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.result_i_tmp_6(result_i_tmp_6),
	.result_i_tmp_5(result_i_tmp_5),
	.result_i_tmp_4(result_i_tmp_4),
	.result_i_tmp_3(result_i_tmp_3),
	.result_i_tmp_2(result_i_tmp_2),
	.result_i_tmp_1(result_i_tmp_1),
	.result_i_tmp_0(result_i_tmp_0),
	.clock(clock));

endmodule

module IFFT_add_sub_8gj_5 (
	clken,
	pipeline_dffe_11,
	pipeline_dffe_15,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	result_i_tmp_11,
	result_i_tmp_15,
	result_i_tmp_12,
	result_i_tmp_13,
	result_i_tmp_14,
	result_i_tmp_10,
	result_i_tmp_9,
	pipeline_dffe_10,
	result_i_tmp_8,
	pipeline_dffe_9,
	result_i_tmp_7,
	pipeline_dffe_8,
	result_i_tmp_6,
	result_i_tmp_5,
	result_i_tmp_4,
	result_i_tmp_3,
	result_i_tmp_2,
	result_i_tmp_1,
	result_i_tmp_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_11;
output 	pipeline_dffe_15;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	result_i_tmp_11;
input 	result_i_tmp_15;
input 	result_i_tmp_12;
input 	result_i_tmp_13;
input 	result_i_tmp_14;
input 	result_i_tmp_10;
input 	result_i_tmp_9;
output 	pipeline_dffe_10;
input 	result_i_tmp_8;
output 	pipeline_dffe_9;
input 	result_i_tmp_7;
output 	pipeline_dffe_8;
input 	result_i_tmp_6;
input 	result_i_tmp_5;
input 	result_i_tmp_4;
input 	result_i_tmp_3;
input 	result_i_tmp_2;
input 	result_i_tmp_1;
input 	result_i_tmp_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[11] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[15] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[12] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[13] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[14] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[10] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!result_i_tmp_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_da2:cm3|u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl_4 (
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_4_1,
	tdl_arr_5_1,
	tdl_arr_6_1,
	data_in,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_4_1;
output 	tdl_arr_5_1;
output 	tdl_arr_6_1;
input 	[7:0] data_in;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][3]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;


dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_5 (
	global_clock_enable,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_4_1,
	tdl_arr_5_1,
	tdl_arr_6_1,
	data_in,
	tdl_arr_2_1,
	tdl_arr_1_1,
	tdl_arr_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	tdl_arr_3_1;
output 	tdl_arr_7_1;
output 	tdl_arr_4_1;
output 	tdl_arr_5_1;
output 	tdl_arr_6_1;
input 	[7:0] data_in;
output 	tdl_arr_2_1;
output 	tdl_arr_1_1;
output 	tdl_arr_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][3]~q ;
wire \tdl_arr[0][7]~q ;
wire \tdl_arr[0][4]~q ;
wire \tdl_arr[0][5]~q ;
wire \tdl_arr[0][6]~q ;
wire \tdl_arr[0][2]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[0][0]~q ;


dffeas \tdl_arr[1][3] (
	.clk(clk),
	.d(\tdl_arr[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_3_1),
	.prn(vcc));
defparam \tdl_arr[1][3] .is_wysiwyg = "true";
defparam \tdl_arr[1][3] .power_up = "low";

dffeas \tdl_arr[1][7] (
	.clk(clk),
	.d(\tdl_arr[0][7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_7_1),
	.prn(vcc));
defparam \tdl_arr[1][7] .is_wysiwyg = "true";
defparam \tdl_arr[1][7] .power_up = "low";

dffeas \tdl_arr[1][4] (
	.clk(clk),
	.d(\tdl_arr[0][4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4_1),
	.prn(vcc));
defparam \tdl_arr[1][4] .is_wysiwyg = "true";
defparam \tdl_arr[1][4] .power_up = "low";

dffeas \tdl_arr[1][5] (
	.clk(clk),
	.d(\tdl_arr[0][5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5_1),
	.prn(vcc));
defparam \tdl_arr[1][5] .is_wysiwyg = "true";
defparam \tdl_arr[1][5] .power_up = "low";

dffeas \tdl_arr[1][6] (
	.clk(clk),
	.d(\tdl_arr[0][6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6_1),
	.prn(vcc));
defparam \tdl_arr[1][6] .is_wysiwyg = "true";
defparam \tdl_arr[1][6] .power_up = "low";

dffeas \tdl_arr[1][2] (
	.clk(clk),
	.d(\tdl_arr[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_2_1),
	.prn(vcc));
defparam \tdl_arr[1][2] .is_wysiwyg = "true";
defparam \tdl_arr[1][2] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_1),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_1),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[0][3] (
	.clk(clk),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][3]~q ),
	.prn(vcc));
defparam \tdl_arr[0][3] .is_wysiwyg = "true";
defparam \tdl_arr[0][3] .power_up = "low";

dffeas \tdl_arr[0][7] (
	.clk(clk),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][7]~q ),
	.prn(vcc));
defparam \tdl_arr[0][7] .is_wysiwyg = "true";
defparam \tdl_arr[0][7] .power_up = "low";

dffeas \tdl_arr[0][4] (
	.clk(clk),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][4]~q ),
	.prn(vcc));
defparam \tdl_arr[0][4] .is_wysiwyg = "true";
defparam \tdl_arr[0][4] .power_up = "low";

dffeas \tdl_arr[0][5] (
	.clk(clk),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][5]~q ),
	.prn(vcc));
defparam \tdl_arr[0][5] .is_wysiwyg = "true";
defparam \tdl_arr[0][5] .power_up = "low";

dffeas \tdl_arr[0][6] (
	.clk(clk),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][6]~q ),
	.prn(vcc));
defparam \tdl_arr[0][6] .is_wysiwyg = "true";
defparam \tdl_arr[0][6] .power_up = "low";

dffeas \tdl_arr[0][2] (
	.clk(clk),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][2]~q ),
	.prn(vcc));
defparam \tdl_arr[0][2] .is_wysiwyg = "true";
defparam \tdl_arr[0][2] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

endmodule

module IFFT_asj_fft_bfp_i (
	r_array_out_2_2,
	r_array_out_2_0,
	i_array_out_2_3,
	i_array_out_2_1,
	r_array_out_3_0,
	r_array_out_3_2,
	i_array_out_3_1,
	i_array_out_3_3,
	r_array_out_4_2,
	r_array_out_4_0,
	i_array_out_4_3,
	i_array_out_4_1,
	r_array_out_5_2,
	r_array_out_5_0,
	i_array_out_5_3,
	i_array_out_5_1,
	r_array_out_2_3,
	r_array_out_2_1,
	i_array_out_2_2,
	i_array_out_2_0,
	r_array_out_3_3,
	r_array_out_3_1,
	i_array_out_3_0,
	i_array_out_3_2,
	r_array_out_4_3,
	r_array_out_4_1,
	i_array_out_4_2,
	i_array_out_4_0,
	i_array_out_5_2,
	i_array_out_5_0,
	r_array_out_5_3,
	r_array_out_5_1,
	r_array_out_1_0,
	r_array_out_1_2,
	i_array_out_1_3,
	i_array_out_1_1,
	r_array_out_1_3,
	r_array_out_1_1,
	i_array_out_1_2,
	i_array_out_1_0,
	r_array_out_0_2,
	r_array_out_0_0,
	i_array_out_0_1,
	i_array_out_0_3,
	r_array_out_0_3,
	r_array_out_0_1,
	i_array_out_0_2,
	i_array_out_0_0,
	global_clock_enable,
	slb_last_0,
	slb_last_1,
	slb_last_2,
	r_array_out_6_1,
	r_array_out_6_3,
	r_array_out_6_0,
	r_array_out_6_2,
	r_array_out_7_1,
	r_array_out_7_3,
	r_array_out_7_0,
	r_array_out_7_2,
	i_array_out_7_1,
	i_array_out_7_3,
	i_array_out_7_0,
	i_array_out_7_2,
	i_array_out_6_1,
	i_array_out_6_3,
	i_array_out_6_0,
	i_array_out_6_2,
	ram_in_reg_6_1,
	ram_in_reg_5_1,
	ram_in_reg_2_1,
	ram_in_reg_3_1,
	ram_in_reg_4_1,
	ram_in_reg_6_3,
	ram_in_reg_5_3,
	ram_in_reg_2_3,
	ram_in_reg_3_3,
	ram_in_reg_4_3,
	ram_in_reg_6_0,
	ram_in_reg_5_0,
	ram_in_reg_2_0,
	ram_in_reg_3_0,
	ram_in_reg_4_0,
	ram_in_reg_6_2,
	ram_in_reg_5_2,
	ram_in_reg_2_2,
	ram_in_reg_3_2,
	ram_in_reg_4_2,
	ram_in_reg_7_1,
	ram_in_reg_7_3,
	ram_in_reg_7_0,
	ram_in_reg_7_2,
	ram_in_reg_7_5,
	ram_in_reg_6_5,
	ram_in_reg_3_5,
	ram_in_reg_4_5,
	ram_in_reg_5_5,
	ram_in_reg_7_7,
	ram_in_reg_6_7,
	ram_in_reg_3_7,
	ram_in_reg_4_7,
	ram_in_reg_5_7,
	ram_in_reg_7_4,
	ram_in_reg_6_4,
	ram_in_reg_3_4,
	ram_in_reg_4_4,
	ram_in_reg_5_4,
	ram_in_reg_7_6,
	ram_in_reg_6_6,
	ram_in_reg_3_6,
	ram_in_reg_4_6,
	ram_in_reg_5_6,
	ram_in_reg_2_5,
	ram_in_reg_2_7,
	ram_in_reg_2_4,
	ram_in_reg_2_6,
	ram_in_reg_0_2,
	ram_in_reg_1_2,
	ram_in_reg_0_0,
	ram_in_reg_1_0,
	ram_in_reg_0_7,
	ram_in_reg_1_7,
	ram_in_reg_0_5,
	ram_in_reg_1_5,
	ram_in_reg_0_3,
	ram_in_reg_1_3,
	ram_in_reg_0_1,
	ram_in_reg_1_1,
	ram_in_reg_0_6,
	ram_in_reg_1_6,
	ram_in_reg_0_4,
	ram_in_reg_1_4,
	clk)/* synthesis synthesis_greybox=1 */;
output 	r_array_out_2_2;
output 	r_array_out_2_0;
output 	i_array_out_2_3;
output 	i_array_out_2_1;
output 	r_array_out_3_0;
output 	r_array_out_3_2;
output 	i_array_out_3_1;
output 	i_array_out_3_3;
output 	r_array_out_4_2;
output 	r_array_out_4_0;
output 	i_array_out_4_3;
output 	i_array_out_4_1;
output 	r_array_out_5_2;
output 	r_array_out_5_0;
output 	i_array_out_5_3;
output 	i_array_out_5_1;
output 	r_array_out_2_3;
output 	r_array_out_2_1;
output 	i_array_out_2_2;
output 	i_array_out_2_0;
output 	r_array_out_3_3;
output 	r_array_out_3_1;
output 	i_array_out_3_0;
output 	i_array_out_3_2;
output 	r_array_out_4_3;
output 	r_array_out_4_1;
output 	i_array_out_4_2;
output 	i_array_out_4_0;
output 	i_array_out_5_2;
output 	i_array_out_5_0;
output 	r_array_out_5_3;
output 	r_array_out_5_1;
output 	r_array_out_1_0;
output 	r_array_out_1_2;
output 	i_array_out_1_3;
output 	i_array_out_1_1;
output 	r_array_out_1_3;
output 	r_array_out_1_1;
output 	i_array_out_1_2;
output 	i_array_out_1_0;
output 	r_array_out_0_2;
output 	r_array_out_0_0;
output 	i_array_out_0_1;
output 	i_array_out_0_3;
output 	r_array_out_0_3;
output 	r_array_out_0_1;
output 	i_array_out_0_2;
output 	i_array_out_0_0;
input 	global_clock_enable;
input 	slb_last_0;
input 	slb_last_1;
input 	slb_last_2;
output 	r_array_out_6_1;
output 	r_array_out_6_3;
output 	r_array_out_6_0;
output 	r_array_out_6_2;
output 	r_array_out_7_1;
output 	r_array_out_7_3;
output 	r_array_out_7_0;
output 	r_array_out_7_2;
output 	i_array_out_7_1;
output 	i_array_out_7_3;
output 	i_array_out_7_0;
output 	i_array_out_7_2;
output 	i_array_out_6_1;
output 	i_array_out_6_3;
output 	i_array_out_6_0;
output 	i_array_out_6_2;
input 	ram_in_reg_6_1;
input 	ram_in_reg_5_1;
input 	ram_in_reg_2_1;
input 	ram_in_reg_3_1;
input 	ram_in_reg_4_1;
input 	ram_in_reg_6_3;
input 	ram_in_reg_5_3;
input 	ram_in_reg_2_3;
input 	ram_in_reg_3_3;
input 	ram_in_reg_4_3;
input 	ram_in_reg_6_0;
input 	ram_in_reg_5_0;
input 	ram_in_reg_2_0;
input 	ram_in_reg_3_0;
input 	ram_in_reg_4_0;
input 	ram_in_reg_6_2;
input 	ram_in_reg_5_2;
input 	ram_in_reg_2_2;
input 	ram_in_reg_3_2;
input 	ram_in_reg_4_2;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_0;
input 	ram_in_reg_7_2;
input 	ram_in_reg_7_5;
input 	ram_in_reg_6_5;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_5;
input 	ram_in_reg_7_7;
input 	ram_in_reg_6_7;
input 	ram_in_reg_3_7;
input 	ram_in_reg_4_7;
input 	ram_in_reg_5_7;
input 	ram_in_reg_7_4;
input 	ram_in_reg_6_4;
input 	ram_in_reg_3_4;
input 	ram_in_reg_4_4;
input 	ram_in_reg_5_4;
input 	ram_in_reg_7_6;
input 	ram_in_reg_6_6;
input 	ram_in_reg_3_6;
input 	ram_in_reg_4_6;
input 	ram_in_reg_5_6;
input 	ram_in_reg_2_5;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_4;
input 	ram_in_reg_2_6;
input 	ram_in_reg_0_2;
input 	ram_in_reg_1_2;
input 	ram_in_reg_0_0;
input 	ram_in_reg_1_0;
input 	ram_in_reg_0_7;
input 	ram_in_reg_1_7;
input 	ram_in_reg_0_5;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_3;
input 	ram_in_reg_1_3;
input 	ram_in_reg_0_1;
input 	ram_in_reg_1_1;
input 	ram_in_reg_0_6;
input 	ram_in_reg_1_6;
input 	ram_in_reg_0_4;
input 	ram_in_reg_1_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux16~3_combout ;
wire \Mux16~4_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux56~3_combout ;
wire \Mux56~4_combout ;
wire \Mux40~3_combout ;
wire \Mux40~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Mux40~5_combout ;
wire \Mux40~6_combout ;
wire \Mux56~5_combout ;
wire \Mux56~6_combout ;
wire \Mux19~0_combout ;
wire \Mux3~0_combout ;
wire \Mux59~0_combout ;
wire \Mux43~0_combout ;
wire \Mux18~0_combout ;
wire \Mux2~0_combout ;
wire \Mux58~0_combout ;
wire \Mux42~0_combout ;
wire \Mux24~3_combout ;
wire \Mux24~4_combout ;
wire \Mux8~3_combout ;
wire \Mux8~4_combout ;
wire \Mux48~3_combout ;
wire \Mux48~4_combout ;
wire \Mux32~3_combout ;
wire \Mux32~4_combout ;
wire \Mux24~5_combout ;
wire \Mux24~6_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \Mux32~5_combout ;
wire \Mux32~6_combout ;
wire \Mux48~5_combout ;
wire \Mux48~6_combout ;
wire \Mux27~0_combout ;
wire \Mux11~0_combout ;
wire \Mux51~0_combout ;
wire \Mux35~0_combout ;
wire \Mux50~0_combout ;
wire \Mux34~0_combout ;
wire \Mux26~0_combout ;
wire \Mux10~0_combout ;
wire \i_array_out[0][6]~1_combout ;
wire \Mux8~0_combout ;
wire \i_array_out[0][6]~0_combout ;
wire \Mux9~0_combout ;
wire \Mux24~0_combout ;
wire \Mux25~0_combout ;
wire \Mux0~0_combout ;
wire \Mux1~0_combout ;
wire \Mux16~0_combout ;
wire \Mux17~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \Mux24~1_combout ;
wire \Mux24~2_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux16~1_combout ;
wire \Mux16~2_combout ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \Mux40~2_combout ;
wire \Mux41~0_combout ;
wire \Mux56~2_combout ;
wire \Mux57~0_combout ;
wire \Mux32~2_combout ;
wire \Mux33~0_combout ;
wire \Mux48~2_combout ;
wire \Mux49~0_combout ;


dffeas \r_array_out[2][2] (
	.clk(clk),
	.d(\Mux16~3_combout ),
	.asdata(\Mux16~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_2_2),
	.prn(vcc));
defparam \r_array_out[2][2] .is_wysiwyg = "true";
defparam \r_array_out[2][2] .power_up = "low";

dffeas \r_array_out[0][2] (
	.clk(clk),
	.d(\Mux0~3_combout ),
	.asdata(\Mux0~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_2_0),
	.prn(vcc));
defparam \r_array_out[0][2] .is_wysiwyg = "true";
defparam \r_array_out[0][2] .power_up = "low";

dffeas \i_array_out[3][2] (
	.clk(clk),
	.d(\Mux56~3_combout ),
	.asdata(\Mux56~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_2_3),
	.prn(vcc));
defparam \i_array_out[3][2] .is_wysiwyg = "true";
defparam \i_array_out[3][2] .power_up = "low";

dffeas \i_array_out[1][2] (
	.clk(clk),
	.d(\Mux40~3_combout ),
	.asdata(\Mux40~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_2_1),
	.prn(vcc));
defparam \i_array_out[1][2] .is_wysiwyg = "true";
defparam \i_array_out[1][2] .power_up = "low";

dffeas \r_array_out[0][3] (
	.clk(clk),
	.d(\Mux0~5_combout ),
	.asdata(\Mux0~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_3_0),
	.prn(vcc));
defparam \r_array_out[0][3] .is_wysiwyg = "true";
defparam \r_array_out[0][3] .power_up = "low";

dffeas \r_array_out[2][3] (
	.clk(clk),
	.d(\Mux16~5_combout ),
	.asdata(\Mux16~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_3_2),
	.prn(vcc));
defparam \r_array_out[2][3] .is_wysiwyg = "true";
defparam \r_array_out[2][3] .power_up = "low";

dffeas \i_array_out[1][3] (
	.clk(clk),
	.d(\Mux40~5_combout ),
	.asdata(\Mux40~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_3_1),
	.prn(vcc));
defparam \i_array_out[1][3] .is_wysiwyg = "true";
defparam \i_array_out[1][3] .power_up = "low";

dffeas \i_array_out[3][3] (
	.clk(clk),
	.d(\Mux56~5_combout ),
	.asdata(\Mux56~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_3_3),
	.prn(vcc));
defparam \i_array_out[3][3] .is_wysiwyg = "true";
defparam \i_array_out[3][3] .power_up = "low";

dffeas \r_array_out[2][4] (
	.clk(clk),
	.d(\Mux19~0_combout ),
	.asdata(ram_in_reg_0_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_4_2),
	.prn(vcc));
defparam \r_array_out[2][4] .is_wysiwyg = "true";
defparam \r_array_out[2][4] .power_up = "low";

dffeas \r_array_out[0][4] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(ram_in_reg_0_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_4_0),
	.prn(vcc));
defparam \r_array_out[0][4] .is_wysiwyg = "true";
defparam \r_array_out[0][4] .power_up = "low";

dffeas \i_array_out[3][4] (
	.clk(clk),
	.d(\Mux59~0_combout ),
	.asdata(ram_in_reg_0_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_4_3),
	.prn(vcc));
defparam \i_array_out[3][4] .is_wysiwyg = "true";
defparam \i_array_out[3][4] .power_up = "low";

dffeas \i_array_out[1][4] (
	.clk(clk),
	.d(\Mux43~0_combout ),
	.asdata(ram_in_reg_0_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_4_1),
	.prn(vcc));
defparam \i_array_out[1][4] .is_wysiwyg = "true";
defparam \i_array_out[1][4] .power_up = "low";

dffeas \r_array_out[2][5] (
	.clk(clk),
	.d(\Mux18~0_combout ),
	.asdata(ram_in_reg_1_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_5_2),
	.prn(vcc));
defparam \r_array_out[2][5] .is_wysiwyg = "true";
defparam \r_array_out[2][5] .power_up = "low";

dffeas \r_array_out[0][5] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(ram_in_reg_1_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_5_0),
	.prn(vcc));
defparam \r_array_out[0][5] .is_wysiwyg = "true";
defparam \r_array_out[0][5] .power_up = "low";

dffeas \i_array_out[3][5] (
	.clk(clk),
	.d(\Mux58~0_combout ),
	.asdata(ram_in_reg_1_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_5_3),
	.prn(vcc));
defparam \i_array_out[3][5] .is_wysiwyg = "true";
defparam \i_array_out[3][5] .power_up = "low";

dffeas \i_array_out[1][5] (
	.clk(clk),
	.d(\Mux42~0_combout ),
	.asdata(ram_in_reg_1_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_5_1),
	.prn(vcc));
defparam \i_array_out[1][5] .is_wysiwyg = "true";
defparam \i_array_out[1][5] .power_up = "low";

dffeas \r_array_out[3][2] (
	.clk(clk),
	.d(\Mux24~3_combout ),
	.asdata(\Mux24~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_2_3),
	.prn(vcc));
defparam \r_array_out[3][2] .is_wysiwyg = "true";
defparam \r_array_out[3][2] .power_up = "low";

dffeas \r_array_out[1][2] (
	.clk(clk),
	.d(\Mux8~3_combout ),
	.asdata(\Mux8~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_2_1),
	.prn(vcc));
defparam \r_array_out[1][2] .is_wysiwyg = "true";
defparam \r_array_out[1][2] .power_up = "low";

dffeas \i_array_out[2][2] (
	.clk(clk),
	.d(\Mux48~3_combout ),
	.asdata(\Mux48~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_2_2),
	.prn(vcc));
defparam \i_array_out[2][2] .is_wysiwyg = "true";
defparam \i_array_out[2][2] .power_up = "low";

dffeas \i_array_out[0][2] (
	.clk(clk),
	.d(\Mux32~3_combout ),
	.asdata(\Mux32~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_2_0),
	.prn(vcc));
defparam \i_array_out[0][2] .is_wysiwyg = "true";
defparam \i_array_out[0][2] .power_up = "low";

dffeas \r_array_out[3][3] (
	.clk(clk),
	.d(\Mux24~5_combout ),
	.asdata(\Mux24~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_3_3),
	.prn(vcc));
defparam \r_array_out[3][3] .is_wysiwyg = "true";
defparam \r_array_out[3][3] .power_up = "low";

dffeas \r_array_out[1][3] (
	.clk(clk),
	.d(\Mux8~5_combout ),
	.asdata(\Mux8~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(r_array_out_3_1),
	.prn(vcc));
defparam \r_array_out[1][3] .is_wysiwyg = "true";
defparam \r_array_out[1][3] .power_up = "low";

dffeas \i_array_out[0][3] (
	.clk(clk),
	.d(\Mux32~5_combout ),
	.asdata(\Mux32~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_3_0),
	.prn(vcc));
defparam \i_array_out[0][3] .is_wysiwyg = "true";
defparam \i_array_out[0][3] .power_up = "low";

dffeas \i_array_out[2][3] (
	.clk(clk),
	.d(\Mux48~5_combout ),
	.asdata(\Mux48~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(slb_last_2),
	.sload(!slb_last_1),
	.ena(!global_clock_enable),
	.q(i_array_out_3_2),
	.prn(vcc));
defparam \i_array_out[2][3] .is_wysiwyg = "true";
defparam \i_array_out[2][3] .power_up = "low";

dffeas \r_array_out[3][4] (
	.clk(clk),
	.d(\Mux27~0_combout ),
	.asdata(ram_in_reg_0_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_4_3),
	.prn(vcc));
defparam \r_array_out[3][4] .is_wysiwyg = "true";
defparam \r_array_out[3][4] .power_up = "low";

dffeas \r_array_out[1][4] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(ram_in_reg_0_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_4_1),
	.prn(vcc));
defparam \r_array_out[1][4] .is_wysiwyg = "true";
defparam \r_array_out[1][4] .power_up = "low";

dffeas \i_array_out[2][4] (
	.clk(clk),
	.d(\Mux51~0_combout ),
	.asdata(ram_in_reg_0_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_4_2),
	.prn(vcc));
defparam \i_array_out[2][4] .is_wysiwyg = "true";
defparam \i_array_out[2][4] .power_up = "low";

dffeas \i_array_out[0][4] (
	.clk(clk),
	.d(\Mux35~0_combout ),
	.asdata(ram_in_reg_0_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_4_0),
	.prn(vcc));
defparam \i_array_out[0][4] .is_wysiwyg = "true";
defparam \i_array_out[0][4] .power_up = "low";

dffeas \i_array_out[2][5] (
	.clk(clk),
	.d(\Mux50~0_combout ),
	.asdata(ram_in_reg_1_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_5_2),
	.prn(vcc));
defparam \i_array_out[2][5] .is_wysiwyg = "true";
defparam \i_array_out[2][5] .power_up = "low";

dffeas \i_array_out[0][5] (
	.clk(clk),
	.d(\Mux34~0_combout ),
	.asdata(ram_in_reg_1_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(i_array_out_5_0),
	.prn(vcc));
defparam \i_array_out[0][5] .is_wysiwyg = "true";
defparam \i_array_out[0][5] .power_up = "low";

dffeas \r_array_out[3][5] (
	.clk(clk),
	.d(\Mux26~0_combout ),
	.asdata(ram_in_reg_1_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_5_3),
	.prn(vcc));
defparam \r_array_out[3][5] .is_wysiwyg = "true";
defparam \r_array_out[3][5] .power_up = "low";

dffeas \r_array_out[1][5] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(ram_in_reg_1_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(slb_last_2),
	.ena(!global_clock_enable),
	.q(r_array_out_5_1),
	.prn(vcc));
defparam \r_array_out[1][5] .is_wysiwyg = "true";
defparam \r_array_out[1][5] .power_up = "low";

dffeas \r_array_out[0][1] (
	.clk(clk),
	.d(\Mux0~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_1_0),
	.prn(vcc));
defparam \r_array_out[0][1] .is_wysiwyg = "true";
defparam \r_array_out[0][1] .power_up = "low";

dffeas \r_array_out[2][1] (
	.clk(clk),
	.d(\Mux16~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_1_2),
	.prn(vcc));
defparam \r_array_out[2][1] .is_wysiwyg = "true";
defparam \r_array_out[2][1] .power_up = "low";

dffeas \i_array_out[3][1] (
	.clk(clk),
	.d(\Mux56~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_1_3),
	.prn(vcc));
defparam \i_array_out[3][1] .is_wysiwyg = "true";
defparam \i_array_out[3][1] .power_up = "low";

dffeas \i_array_out[1][1] (
	.clk(clk),
	.d(\Mux40~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_1_1),
	.prn(vcc));
defparam \i_array_out[1][1] .is_wysiwyg = "true";
defparam \i_array_out[1][1] .power_up = "low";

dffeas \r_array_out[3][1] (
	.clk(clk),
	.d(\Mux24~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_1_3),
	.prn(vcc));
defparam \r_array_out[3][1] .is_wysiwyg = "true";
defparam \r_array_out[3][1] .power_up = "low";

dffeas \r_array_out[1][1] (
	.clk(clk),
	.d(\Mux8~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_1_1),
	.prn(vcc));
defparam \r_array_out[1][1] .is_wysiwyg = "true";
defparam \r_array_out[1][1] .power_up = "low";

dffeas \i_array_out[2][1] (
	.clk(clk),
	.d(\Mux48~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_1_2),
	.prn(vcc));
defparam \i_array_out[2][1] .is_wysiwyg = "true";
defparam \i_array_out[2][1] .power_up = "low";

dffeas \i_array_out[0][1] (
	.clk(clk),
	.d(\Mux32~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_1_0),
	.prn(vcc));
defparam \i_array_out[0][1] .is_wysiwyg = "true";
defparam \i_array_out[0][1] .power_up = "low";

dffeas \r_array_out[2][0] (
	.clk(clk),
	.d(\Mux16~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_0_2),
	.prn(vcc));
defparam \r_array_out[2][0] .is_wysiwyg = "true";
defparam \r_array_out[2][0] .power_up = "low";

dffeas \r_array_out[0][0] (
	.clk(clk),
	.d(\Mux0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_0_0),
	.prn(vcc));
defparam \r_array_out[0][0] .is_wysiwyg = "true";
defparam \r_array_out[0][0] .power_up = "low";

dffeas \i_array_out[1][0] (
	.clk(clk),
	.d(\Mux40~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_0_1),
	.prn(vcc));
defparam \i_array_out[1][0] .is_wysiwyg = "true";
defparam \i_array_out[1][0] .power_up = "low";

dffeas \i_array_out[3][0] (
	.clk(clk),
	.d(\Mux56~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_0_3),
	.prn(vcc));
defparam \i_array_out[3][0] .is_wysiwyg = "true";
defparam \i_array_out[3][0] .power_up = "low";

dffeas \r_array_out[3][0] (
	.clk(clk),
	.d(\Mux24~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_0_3),
	.prn(vcc));
defparam \r_array_out[3][0] .is_wysiwyg = "true";
defparam \r_array_out[3][0] .power_up = "low";

dffeas \r_array_out[1][0] (
	.clk(clk),
	.d(\Mux8~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_0_1),
	.prn(vcc));
defparam \r_array_out[1][0] .is_wysiwyg = "true";
defparam \r_array_out[1][0] .power_up = "low";

dffeas \i_array_out[2][0] (
	.clk(clk),
	.d(\Mux48~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_0_2),
	.prn(vcc));
defparam \i_array_out[2][0] .is_wysiwyg = "true";
defparam \i_array_out[2][0] .power_up = "low";

dffeas \i_array_out[0][0] (
	.clk(clk),
	.d(\Mux32~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\i_array_out[0][6]~1_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_0_0),
	.prn(vcc));
defparam \i_array_out[0][0] .is_wysiwyg = "true";
defparam \i_array_out[0][0] .power_up = "low";

dffeas \r_array_out[1][6] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_6_1),
	.prn(vcc));
defparam \r_array_out[1][6] .is_wysiwyg = "true";
defparam \r_array_out[1][6] .power_up = "low";

dffeas \r_array_out[3][6] (
	.clk(clk),
	.d(\Mux25~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_6_3),
	.prn(vcc));
defparam \r_array_out[3][6] .is_wysiwyg = "true";
defparam \r_array_out[3][6] .power_up = "low";

dffeas \r_array_out[0][6] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_6_0),
	.prn(vcc));
defparam \r_array_out[0][6] .is_wysiwyg = "true";
defparam \r_array_out[0][6] .power_up = "low";

dffeas \r_array_out[2][6] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_6_2),
	.prn(vcc));
defparam \r_array_out[2][6] .is_wysiwyg = "true";
defparam \r_array_out[2][6] .power_up = "low";

dffeas \r_array_out[1][7] (
	.clk(clk),
	.d(\Mux8~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_7_1),
	.prn(vcc));
defparam \r_array_out[1][7] .is_wysiwyg = "true";
defparam \r_array_out[1][7] .power_up = "low";

dffeas \r_array_out[3][7] (
	.clk(clk),
	.d(\Mux24~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_7_3),
	.prn(vcc));
defparam \r_array_out[3][7] .is_wysiwyg = "true";
defparam \r_array_out[3][7] .power_up = "low";

dffeas \r_array_out[0][7] (
	.clk(clk),
	.d(\Mux0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_7_0),
	.prn(vcc));
defparam \r_array_out[0][7] .is_wysiwyg = "true";
defparam \r_array_out[0][7] .power_up = "low";

dffeas \r_array_out[2][7] (
	.clk(clk),
	.d(\Mux16~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(r_array_out_7_2),
	.prn(vcc));
defparam \r_array_out[2][7] .is_wysiwyg = "true";
defparam \r_array_out[2][7] .power_up = "low";

dffeas \i_array_out[1][7] (
	.clk(clk),
	.d(\Mux40~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_7_1),
	.prn(vcc));
defparam \i_array_out[1][7] .is_wysiwyg = "true";
defparam \i_array_out[1][7] .power_up = "low";

dffeas \i_array_out[3][7] (
	.clk(clk),
	.d(\Mux56~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_7_3),
	.prn(vcc));
defparam \i_array_out[3][7] .is_wysiwyg = "true";
defparam \i_array_out[3][7] .power_up = "low";

dffeas \i_array_out[0][7] (
	.clk(clk),
	.d(\Mux32~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_7_0),
	.prn(vcc));
defparam \i_array_out[0][7] .is_wysiwyg = "true";
defparam \i_array_out[0][7] .power_up = "low";

dffeas \i_array_out[2][7] (
	.clk(clk),
	.d(\Mux48~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_7_2),
	.prn(vcc));
defparam \i_array_out[2][7] .is_wysiwyg = "true";
defparam \i_array_out[2][7] .power_up = "low";

dffeas \i_array_out[1][6] (
	.clk(clk),
	.d(\Mux41~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_6_1),
	.prn(vcc));
defparam \i_array_out[1][6] .is_wysiwyg = "true";
defparam \i_array_out[1][6] .power_up = "low";

dffeas \i_array_out[3][6] (
	.clk(clk),
	.d(\Mux57~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_6_3),
	.prn(vcc));
defparam \i_array_out[3][6] .is_wysiwyg = "true";
defparam \i_array_out[3][6] .power_up = "low";

dffeas \i_array_out[0][6] (
	.clk(clk),
	.d(\Mux33~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_6_0),
	.prn(vcc));
defparam \i_array_out[0][6] .is_wysiwyg = "true";
defparam \i_array_out[0][6] .power_up = "low";

dffeas \i_array_out[2][6] (
	.clk(clk),
	.d(\Mux49~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(i_array_out_6_2),
	.prn(vcc));
defparam \i_array_out[2][6] .is_wysiwyg = "true";
defparam \i_array_out[2][6] .power_up = "low";

cyclonev_lcell_comb \Mux16~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~3 .extended_lut = "off";
defparam \Mux16~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux16~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_2),
	.datac(!ram_in_reg_1_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~4 .extended_lut = "off";
defparam \Mux16~4 .lut_mask = 64'h2727272727272727;
defparam \Mux16~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~3 .extended_lut = "off";
defparam \Mux0~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux0~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_0),
	.datac(!ram_in_reg_1_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~4 .extended_lut = "off";
defparam \Mux0~4 .lut_mask = 64'h2727272727272727;
defparam \Mux0~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~3 .extended_lut = "off";
defparam \Mux56~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux56~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_7),
	.datac(!ram_in_reg_1_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~4 .extended_lut = "off";
defparam \Mux56~4 .lut_mask = 64'h2727272727272727;
defparam \Mux56~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~3 .extended_lut = "off";
defparam \Mux40~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux40~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_5),
	.datac(!ram_in_reg_1_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~4 .extended_lut = "off";
defparam \Mux40~4 .lut_mask = 64'h2727272727272727;
defparam \Mux40~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_0),
	.datac(!ram_in_reg_0_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~5 .extended_lut = "off";
defparam \Mux0~5 .lut_mask = 64'h2727272727272727;
defparam \Mux0~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_0),
	.datac(!ram_in_reg_3_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~6 .extended_lut = "off";
defparam \Mux0~6 .lut_mask = 64'h2727272727272727;
defparam \Mux0~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_2),
	.datac(!ram_in_reg_0_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~5 .extended_lut = "off";
defparam \Mux16~5 .lut_mask = 64'h2727272727272727;
defparam \Mux16~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_2),
	.datac(!ram_in_reg_3_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~6 .extended_lut = "off";
defparam \Mux16~6 .lut_mask = 64'h2727272727272727;
defparam \Mux16~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_5),
	.datac(!ram_in_reg_0_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~5 .extended_lut = "off";
defparam \Mux40~5 .lut_mask = 64'h2727272727272727;
defparam \Mux40~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_5),
	.datac(!ram_in_reg_2_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~6 .extended_lut = "off";
defparam \Mux40~6 .lut_mask = 64'h2727272727272727;
defparam \Mux40~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_7),
	.datac(!ram_in_reg_0_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~5 .extended_lut = "off";
defparam \Mux56~5 .lut_mask = 64'h2727272727272727;
defparam \Mux56~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_7),
	.datac(!ram_in_reg_2_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~6 .extended_lut = "off";
defparam \Mux56~6 .lut_mask = 64'h2727272727272727;
defparam \Mux56~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux19~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_2_2),
	.datad(!ram_in_reg_3_2),
	.datae(!ram_in_reg_4_2),
	.dataf(!ram_in_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux19~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_2_0),
	.datad(!ram_in_reg_3_0),
	.datae(!ram_in_reg_4_0),
	.dataf(!ram_in_reg_1_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux59~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_7),
	.datad(!ram_in_reg_4_7),
	.datae(!ram_in_reg_2_7),
	.dataf(!ram_in_reg_1_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux59~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux59~0 .extended_lut = "off";
defparam \Mux59~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux59~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux43~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_5),
	.datad(!ram_in_reg_4_5),
	.datae(!ram_in_reg_2_5),
	.dataf(!ram_in_reg_1_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux43~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux43~0 .extended_lut = "off";
defparam \Mux43~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux43~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux18~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_5_2),
	.datad(!ram_in_reg_2_2),
	.datae(!ram_in_reg_3_2),
	.dataf(!ram_in_reg_4_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux18~0 .extended_lut = "off";
defparam \Mux18~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux18~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_5_0),
	.datad(!ram_in_reg_2_0),
	.datae(!ram_in_reg_3_0),
	.dataf(!ram_in_reg_4_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux58~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_7),
	.datad(!ram_in_reg_4_7),
	.datae(!ram_in_reg_5_7),
	.dataf(!ram_in_reg_2_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux58~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux58~0 .extended_lut = "off";
defparam \Mux58~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux58~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux42~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_5),
	.datad(!ram_in_reg_4_5),
	.datae(!ram_in_reg_5_5),
	.dataf(!ram_in_reg_2_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux42~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux42~0 .extended_lut = "off";
defparam \Mux42~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux42~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~3 .extended_lut = "off";
defparam \Mux24~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux24~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_3),
	.datac(!ram_in_reg_1_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~4 .extended_lut = "off";
defparam \Mux24~4 .lut_mask = 64'h2727272727272727;
defparam \Mux24~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~3 .extended_lut = "off";
defparam \Mux8~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux8~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_1),
	.datac(!ram_in_reg_1_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~4 .extended_lut = "off";
defparam \Mux8~4 .lut_mask = 64'h2727272727272727;
defparam \Mux8~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~3 .extended_lut = "off";
defparam \Mux48~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux48~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_6),
	.datac(!ram_in_reg_1_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~4 .extended_lut = "off";
defparam \Mux48~4 .lut_mask = 64'h2727272727272727;
defparam \Mux48~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~3 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_0_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~3 .extended_lut = "off";
defparam \Mux32~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux32~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~4 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_4),
	.datac(!ram_in_reg_1_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~4 .extended_lut = "off";
defparam \Mux32~4 .lut_mask = 64'h2727272727272727;
defparam \Mux32~4 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_3),
	.datac(!ram_in_reg_0_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~5 .extended_lut = "off";
defparam \Mux24~5 .lut_mask = 64'h2727272727272727;
defparam \Mux24~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_3),
	.datac(!ram_in_reg_3_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~6 .extended_lut = "off";
defparam \Mux24~6 .lut_mask = 64'h2727272727272727;
defparam \Mux24~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_1),
	.datac(!ram_in_reg_0_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~5 .extended_lut = "off";
defparam \Mux8~5 .lut_mask = 64'h2727272727272727;
defparam \Mux8~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_2_1),
	.datac(!ram_in_reg_3_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~6 .extended_lut = "off";
defparam \Mux8~6 .lut_mask = 64'h2727272727272727;
defparam \Mux8~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_4),
	.datac(!ram_in_reg_0_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~5 .extended_lut = "off";
defparam \Mux32~5 .lut_mask = 64'h2727272727272727;
defparam \Mux32~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_4),
	.datac(!ram_in_reg_2_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~6 .extended_lut = "off";
defparam \Mux32~6 .lut_mask = 64'h2727272727272727;
defparam \Mux32~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~5 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_1_6),
	.datac(!ram_in_reg_0_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~5 .extended_lut = "off";
defparam \Mux48~5 .lut_mask = 64'h2727272727272727;
defparam \Mux48~5 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~6 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_6),
	.datac(!ram_in_reg_2_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~6 .extended_lut = "off";
defparam \Mux48~6 .lut_mask = 64'h2727272727272727;
defparam \Mux48~6 .shared_arith = "off";

cyclonev_lcell_comb \Mux27~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_2_3),
	.datad(!ram_in_reg_3_3),
	.datae(!ram_in_reg_4_3),
	.dataf(!ram_in_reg_1_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux27~0 .extended_lut = "off";
defparam \Mux27~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux27~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_2_1),
	.datad(!ram_in_reg_3_1),
	.datae(!ram_in_reg_4_1),
	.dataf(!ram_in_reg_1_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux51~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_6),
	.datad(!ram_in_reg_4_6),
	.datae(!ram_in_reg_2_6),
	.dataf(!ram_in_reg_1_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux51~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux51~0 .extended_lut = "off";
defparam \Mux51~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux51~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux35~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_4),
	.datad(!ram_in_reg_4_4),
	.datae(!ram_in_reg_2_4),
	.dataf(!ram_in_reg_1_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux35~0 .extended_lut = "off";
defparam \Mux35~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux35~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux50~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_6),
	.datad(!ram_in_reg_4_6),
	.datae(!ram_in_reg_5_6),
	.dataf(!ram_in_reg_2_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux50~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux50~0 .extended_lut = "off";
defparam \Mux50~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux50~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux34~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_3_4),
	.datad(!ram_in_reg_4_4),
	.datae(!ram_in_reg_5_4),
	.dataf(!ram_in_reg_2_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux34~0 .extended_lut = "off";
defparam \Mux34~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux34~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux26~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_5_3),
	.datad(!ram_in_reg_2_3),
	.datae(!ram_in_reg_3_3),
	.dataf(!ram_in_reg_4_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux26~0 .extended_lut = "off";
defparam \Mux26~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux26~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!ram_in_reg_5_1),
	.datad(!ram_in_reg_2_1),
	.datae(!ram_in_reg_3_1),
	.dataf(!ram_in_reg_4_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \i_array_out[0][6]~1 (
	.dataa(!slb_last_1),
	.datab(!slb_last_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_array_out[0][6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_array_out[0][6]~1 .extended_lut = "off";
defparam \i_array_out[0][6]~1 .lut_mask = 64'h7777777777777777;
defparam \i_array_out[0][6]~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_1),
	.datac(!ram_in_reg_4_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h2727272727272727;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \i_array_out[0][6]~0 (
	.dataa(!slb_last_0),
	.datab(!slb_last_1),
	.datac(!slb_last_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_array_out[0][6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_array_out[0][6]~0 .extended_lut = "off";
defparam \i_array_out[0][6]~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \i_array_out[0][6]~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!ram_in_reg_6_1),
	.datab(!ram_in_reg_5_1),
	.datac(!ram_in_reg_2_1),
	.datad(!\Mux8~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_3),
	.datac(!ram_in_reg_4_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~0 .extended_lut = "off";
defparam \Mux24~0 .lut_mask = 64'h2727272727272727;
defparam \Mux24~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux25~0 (
	.dataa(!ram_in_reg_6_3),
	.datab(!ram_in_reg_5_3),
	.datac(!ram_in_reg_2_3),
	.datad(!\Mux24~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "off";
defparam \Mux25~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux25~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_0),
	.datac(!ram_in_reg_4_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h2727272727272727;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!ram_in_reg_6_0),
	.datab(!ram_in_reg_5_0),
	.datac(!ram_in_reg_2_0),
	.datad(!\Mux0~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_2),
	.datac(!ram_in_reg_4_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "off";
defparam \Mux16~0 .lut_mask = 64'h2727272727272727;
defparam \Mux16~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux17~0 (
	.dataa(!ram_in_reg_6_2),
	.datab(!ram_in_reg_5_2),
	.datac(!ram_in_reg_2_2),
	.datad(!\Mux16~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux17~0 .extended_lut = "off";
defparam \Mux17~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux17~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~1 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_5_1),
	.datac(!ram_in_reg_4_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~1 .extended_lut = "off";
defparam \Mux8~1 .lut_mask = 64'h2727272727272727;
defparam \Mux8~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~2 (
	.dataa(!ram_in_reg_7_1),
	.datab(!ram_in_reg_6_1),
	.datac(!ram_in_reg_3_1),
	.datad(!\Mux8~1_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~2 .extended_lut = "off";
defparam \Mux8~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~1 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_5_3),
	.datac(!ram_in_reg_4_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~1 .extended_lut = "off";
defparam \Mux24~1 .lut_mask = 64'h2727272727272727;
defparam \Mux24~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux24~2 (
	.dataa(!ram_in_reg_7_3),
	.datab(!ram_in_reg_6_3),
	.datac(!ram_in_reg_3_3),
	.datad(!\Mux24~1_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux24~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux24~2 .extended_lut = "off";
defparam \Mux24~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux24~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_5_0),
	.datac(!ram_in_reg_4_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'h2727272727272727;
defparam \Mux0~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~2 (
	.dataa(!ram_in_reg_7_0),
	.datab(!ram_in_reg_6_0),
	.datac(!ram_in_reg_3_0),
	.datad(!\Mux0~1_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~2 .extended_lut = "off";
defparam \Mux0~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~1 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_5_2),
	.datac(!ram_in_reg_4_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~1 .extended_lut = "off";
defparam \Mux16~1 .lut_mask = 64'h2727272727272727;
defparam \Mux16~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux16~2 (
	.dataa(!ram_in_reg_7_2),
	.datab(!ram_in_reg_6_2),
	.datac(!ram_in_reg_3_2),
	.datad(!\Mux16~1_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~2 .extended_lut = "off";
defparam \Mux16~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux16~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_4_5),
	.datac(!ram_in_reg_5_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~0 .extended_lut = "off";
defparam \Mux40~0 .lut_mask = 64'h2727272727272727;
defparam \Mux40~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~1 (
	.dataa(!ram_in_reg_7_5),
	.datab(!ram_in_reg_6_5),
	.datac(!ram_in_reg_3_5),
	.datad(!\Mux40~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~1 .extended_lut = "off";
defparam \Mux40~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux40~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_4_7),
	.datac(!ram_in_reg_5_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~0 .extended_lut = "off";
defparam \Mux56~0 .lut_mask = 64'h2727272727272727;
defparam \Mux56~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~1 (
	.dataa(!ram_in_reg_7_7),
	.datab(!ram_in_reg_6_7),
	.datac(!ram_in_reg_3_7),
	.datad(!\Mux56~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~1 .extended_lut = "off";
defparam \Mux56~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux56~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_4_4),
	.datac(!ram_in_reg_5_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~0 .extended_lut = "off";
defparam \Mux32~0 .lut_mask = 64'h2727272727272727;
defparam \Mux32~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~1 (
	.dataa(!ram_in_reg_7_4),
	.datab(!ram_in_reg_6_4),
	.datac(!ram_in_reg_3_4),
	.datad(!\Mux32~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~1 .extended_lut = "off";
defparam \Mux32~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux32~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~0 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_4_6),
	.datac(!ram_in_reg_5_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~0 .extended_lut = "off";
defparam \Mux48~0 .lut_mask = 64'h2727272727272727;
defparam \Mux48~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~1 (
	.dataa(!ram_in_reg_7_6),
	.datab(!ram_in_reg_6_6),
	.datac(!ram_in_reg_3_6),
	.datad(!\Mux48~0_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~1 .extended_lut = "off";
defparam \Mux48~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux48~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux40~2 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_5),
	.datac(!ram_in_reg_4_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux40~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux40~2 .extended_lut = "off";
defparam \Mux40~2 .lut_mask = 64'h2727272727272727;
defparam \Mux40~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux41~0 (
	.dataa(!ram_in_reg_6_5),
	.datab(!ram_in_reg_5_5),
	.datac(!ram_in_reg_2_5),
	.datad(!\Mux40~2_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux41~0 .extended_lut = "off";
defparam \Mux41~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux41~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux56~2 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_7),
	.datac(!ram_in_reg_4_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux56~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux56~2 .extended_lut = "off";
defparam \Mux56~2 .lut_mask = 64'h2727272727272727;
defparam \Mux56~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux57~0 (
	.dataa(!ram_in_reg_6_7),
	.datab(!ram_in_reg_5_7),
	.datac(!ram_in_reg_2_7),
	.datad(!\Mux56~2_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux57~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux57~0 .extended_lut = "off";
defparam \Mux57~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux57~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux32~2 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_4),
	.datac(!ram_in_reg_4_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux32~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux32~2 .extended_lut = "off";
defparam \Mux32~2 .lut_mask = 64'h2727272727272727;
defparam \Mux32~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux33~0 (
	.dataa(!ram_in_reg_6_4),
	.datab(!ram_in_reg_5_4),
	.datac(!ram_in_reg_2_4),
	.datad(!\Mux32~2_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux33~0 .extended_lut = "off";
defparam \Mux33~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux33~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux48~2 (
	.dataa(!slb_last_0),
	.datab(!ram_in_reg_3_6),
	.datac(!ram_in_reg_4_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux48~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux48~2 .extended_lut = "off";
defparam \Mux48~2 .lut_mask = 64'h2727272727272727;
defparam \Mux48~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux49~0 (
	.dataa(!ram_in_reg_6_6),
	.datab(!ram_in_reg_5_6),
	.datac(!ram_in_reg_2_6),
	.datad(!\Mux48~2_combout ),
	.datae(!\i_array_out[0][6]~0_combout ),
	.dataf(!\i_array_out[0][6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux49~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux49~0 .extended_lut = "off";
defparam \Mux49~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux49~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_bfp_o (
	next_block,
	reg_no_twiddle603,
	reg_no_twiddle607,
	reg_no_twiddle617,
	reg_no_twiddle613,
	reg_no_twiddle604,
	reg_no_twiddle614,
	reg_no_twiddle605,
	reg_no_twiddle615,
	reg_no_twiddle606,
	reg_no_twiddle616,
	tdl_arr_9,
	global_clock_enable,
	lut_out_tmp_0,
	lut_out_tmp_1,
	lut_out_tmp_2,
	tdl_arr_3_1,
	tdl_arr_7_1,
	tdl_arr_3_11,
	tdl_arr_7_11,
	tdl_arr_3_12,
	tdl_arr_7_12,
	tdl_arr_3_13,
	tdl_arr_7_13,
	tdl_arr_3_14,
	tdl_arr_7_14,
	tdl_arr_3_15,
	tdl_arr_7_15,
	tdl_arr_4_1,
	tdl_arr_4_11,
	tdl_arr_4_12,
	tdl_arr_4_13,
	tdl_arr_4_14,
	tdl_arr_4_15,
	tdl_arr_5_1,
	tdl_arr_5_11,
	tdl_arr_5_12,
	tdl_arr_5_13,
	tdl_arr_5_14,
	tdl_arr_5_15,
	tdl_arr_6_1,
	tdl_arr_6_11,
	tdl_arr_6_12,
	tdl_arr_6_13,
	tdl_arr_6_14,
	tdl_arr_6_15,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	next_block;
input 	reg_no_twiddle603;
input 	reg_no_twiddle607;
input 	reg_no_twiddle617;
input 	reg_no_twiddle613;
input 	reg_no_twiddle604;
input 	reg_no_twiddle614;
input 	reg_no_twiddle605;
input 	reg_no_twiddle615;
input 	reg_no_twiddle606;
input 	reg_no_twiddle616;
input 	tdl_arr_9;
input 	global_clock_enable;
output 	lut_out_tmp_0;
output 	lut_out_tmp_1;
output 	lut_out_tmp_2;
input 	tdl_arr_3_1;
input 	tdl_arr_7_1;
input 	tdl_arr_3_11;
input 	tdl_arr_7_11;
input 	tdl_arr_3_12;
input 	tdl_arr_7_12;
input 	tdl_arr_3_13;
input 	tdl_arr_7_13;
input 	tdl_arr_3_14;
input 	tdl_arr_7_14;
input 	tdl_arr_3_15;
input 	tdl_arr_7_15;
input 	tdl_arr_4_1;
input 	tdl_arr_4_11;
input 	tdl_arr_4_12;
input 	tdl_arr_4_13;
input 	tdl_arr_4_14;
input 	tdl_arr_4_15;
input 	tdl_arr_5_1;
input 	tdl_arr_5_11;
input 	tdl_arr_5_12;
input 	tdl_arr_5_13;
input 	tdl_arr_5_14;
input 	tdl_arr_5_15;
input 	tdl_arr_6_1;
input 	tdl_arr_6_11;
input 	tdl_arr_6_12;
input 	tdl_arr_6_13;
input 	tdl_arr_6_14;
input 	tdl_arr_6_15;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_blk_float:gen_streaming:gen_disc:delay_next_blk|tdl_arr[0]~q ;
wire \gen_blk_float:gen_streaming:gen_disc:gen_consts_64:delay_next_pass|tdl_arr[6]~q ;
wire \sdetd.IDLE~q ;
wire \Equal0~0_combout ;
wire \sdetd.BLOCK_READY~0_combout ;
wire \sdetd.BLOCK_READY~1_combout ;
wire \sdetd.BLOCK_READY~q ;
wire \sdetd.SLBI~0_combout ;
wire \sdetd.SLBI~q ;
wire \Equal1~0_combout ;
wire \sdetd.DISABLE~0_combout ;
wire \sdetd.DISABLE~q ;
wire \del_np_cnt[2]~0_combout ;
wire \del_np_cnt~1_combout ;
wire \del_np_cnt[0]~q ;
wire \del_np_cnt~5_combout ;
wire \del_np_cnt[1]~q ;
wire \del_np_cnt~4_combout ;
wire \del_np_cnt[2]~q ;
wire \del_np_cnt~3_combout ;
wire \del_np_cnt[3]~q ;
wire \del_np_cnt~2_combout ;
wire \del_np_cnt[4]~q ;
wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \sdetd.ENABLE~q ;
wire \sdetd~8_combout ;
wire \sdetd.GBLK~q ;
wire \gain_lut_8pts~0_combout ;
wire \gain_lut_8pts~1_combout ;
wire \gain_lut_8pts~2_combout ;
wire \gain_lut_8pts~3_combout ;
wire \gain_lut_8pts[0]~q ;
wire \Selector6~0_combout ;
wire \gain_lut_blk[0]~q ;
wire \slb_i[0]~combout ;
wire \gain_lut_8pts~4_combout ;
wire \gain_lut_8pts~5_combout ;
wire \gain_lut_8pts~6_combout ;
wire \gain_lut_8pts~7_combout ;
wire \gain_lut_8pts[1]~q ;
wire \Selector5~0_combout ;
wire \gain_lut_blk[1]~q ;
wire \slb_i[1]~combout ;
wire \gain_lut_8pts~8_combout ;
wire \gain_lut_8pts~9_combout ;
wire \gain_lut_8pts~10_combout ;
wire \gain_lut_8pts~11_combout ;
wire \gain_lut_8pts[2]~q ;
wire \Selector4~0_combout ;
wire \gain_lut_blk[2]~q ;
wire \slb_i[2]~combout ;
wire \gain_lut_8pts~12_combout ;
wire \gain_lut_8pts~13_combout ;
wire \gain_lut_8pts~14_combout ;
wire \gain_lut_8pts~15_combout ;
wire \gain_lut_8pts[3]~q ;
wire \Selector3~0_combout ;
wire \gain_lut_blk[3]~q ;
wire \slb_i[3]~combout ;
wire \lut_out_tmp~0_combout ;
wire \lut_out_tmp[2]~1_combout ;
wire \lut_out_tmp~2_combout ;
wire \lut_out_tmp~3_combout ;


IFFT_asj_fft_tdl_bit_rst_3 \gen_blk_float:gen_streaming:gen_disc:gen_consts_64:delay_next_pass (
	.tdl_arr_6(\gen_blk_float:gen_streaming:gen_disc:gen_consts_64:delay_next_pass|tdl_arr[6]~q ),
	.tdl_arr_9(tdl_arr_9),
	.global_clock_enable(global_clock_enable),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_tdl_bit_rst_2 \gen_blk_float:gen_streaming:gen_disc:delay_next_blk (
	.next_block(next_block),
	.tdl_arr_0(\gen_blk_float:gen_streaming:gen_disc:delay_next_blk|tdl_arr[0]~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk),
	.reset_n(reset_n));

dffeas \lut_out_tmp[0] (
	.clk(clk),
	.d(\lut_out_tmp~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\lut_out_tmp[2]~1_combout ),
	.q(lut_out_tmp_0),
	.prn(vcc));
defparam \lut_out_tmp[0] .is_wysiwyg = "true";
defparam \lut_out_tmp[0] .power_up = "low";

dffeas \lut_out_tmp[1] (
	.clk(clk),
	.d(\lut_out_tmp~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\lut_out_tmp[2]~1_combout ),
	.q(lut_out_tmp_1),
	.prn(vcc));
defparam \lut_out_tmp[1] .is_wysiwyg = "true";
defparam \lut_out_tmp[1] .power_up = "low";

dffeas \lut_out_tmp[2] (
	.clk(clk),
	.d(\lut_out_tmp~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\lut_out_tmp[2]~1_combout ),
	.q(lut_out_tmp_2),
	.prn(vcc));
defparam \lut_out_tmp[2] .is_wysiwyg = "true";
defparam \lut_out_tmp[2] .power_up = "low";

dffeas \sdetd.IDLE (
	.clk(clk),
	.d(reset_n),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sdetd.IDLE~q ),
	.prn(vcc));
defparam \sdetd.IDLE .is_wysiwyg = "true";
defparam \sdetd.IDLE .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\del_np_cnt[4]~q ),
	.datab(!\del_np_cnt[3]~q ),
	.datac(!\del_np_cnt[2]~q ),
	.datad(!\del_np_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \sdetd.BLOCK_READY~0 (
	.dataa(!global_clock_enable),
	.datab(!\sdetd.BLOCK_READY~q ),
	.datac(!\del_np_cnt[0]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdetd.BLOCK_READY~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdetd.BLOCK_READY~0 .extended_lut = "off";
defparam \sdetd.BLOCK_READY~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sdetd.BLOCK_READY~0 .shared_arith = "off";

cyclonev_lcell_comb \sdetd.BLOCK_READY~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\sdetd.ENABLE~q ),
	.datad(!\gen_blk_float:gen_streaming:gen_disc:delay_next_blk|tdl_arr[0]~q ),
	.datae(!\gen_blk_float:gen_streaming:gen_disc:gen_consts_64:delay_next_pass|tdl_arr[6]~q ),
	.dataf(!\sdetd.BLOCK_READY~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdetd.BLOCK_READY~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdetd.BLOCK_READY~1 .extended_lut = "off";
defparam \sdetd.BLOCK_READY~1 .lut_mask = 64'hDFFF1FFFFFFFFFFF;
defparam \sdetd.BLOCK_READY~1 .shared_arith = "off";

dffeas \sdetd.BLOCK_READY (
	.clk(clk),
	.d(\sdetd.BLOCK_READY~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sdetd.BLOCK_READY~q ),
	.prn(vcc));
defparam \sdetd.BLOCK_READY .is_wysiwyg = "true";
defparam \sdetd.BLOCK_READY .power_up = "low";

cyclonev_lcell_comb \sdetd.SLBI~0 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\sdetd.SLBI~q ),
	.datad(!\sdetd.GBLK~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdetd.SLBI~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdetd.SLBI~0 .extended_lut = "off";
defparam \sdetd.SLBI~0 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \sdetd.SLBI~0 .shared_arith = "off";

dffeas \sdetd.SLBI (
	.clk(clk),
	.d(\sdetd.SLBI~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sdetd.SLBI~q ),
	.prn(vcc));
defparam \sdetd.SLBI .is_wysiwyg = "true";
defparam \sdetd.SLBI .power_up = "low";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!\del_np_cnt[4]~q ),
	.datab(!\del_np_cnt[3]~q ),
	.datac(!\del_np_cnt[2]~q ),
	.datad(!\del_np_cnt[1]~q ),
	.datae(!\del_np_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \sdetd.DISABLE~0 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\sdetd.SLBI~q ),
	.datad(!\sdetd.DISABLE~q ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdetd.DISABLE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdetd.DISABLE~0 .extended_lut = "off";
defparam \sdetd.DISABLE~0 .lut_mask = 64'hDFFF1FFFDFFF1FFF;
defparam \sdetd.DISABLE~0 .shared_arith = "off";

dffeas \sdetd.DISABLE (
	.clk(clk),
	.d(\sdetd.DISABLE~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sdetd.DISABLE~q ),
	.prn(vcc));
defparam \sdetd.DISABLE .is_wysiwyg = "true";
defparam \sdetd.DISABLE .power_up = "low";

cyclonev_lcell_comb \del_np_cnt[2]~0 (
	.dataa(!reset_n),
	.datab(!\sdetd.BLOCK_READY~q ),
	.datac(!\sdetd.DISABLE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_np_cnt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_np_cnt[2]~0 .extended_lut = "off";
defparam \del_np_cnt[2]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \del_np_cnt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \del_np_cnt~1 (
	.dataa(!\del_np_cnt[0]~q ),
	.datab(!\del_np_cnt[2]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_np_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_np_cnt~1 .extended_lut = "off";
defparam \del_np_cnt~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \del_np_cnt~1 .shared_arith = "off";

dffeas \del_np_cnt[0] (
	.clk(clk),
	.d(\del_np_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_np_cnt[0]~q ),
	.prn(vcc));
defparam \del_np_cnt[0] .is_wysiwyg = "true";
defparam \del_np_cnt[0] .power_up = "low";

cyclonev_lcell_comb \del_np_cnt~5 (
	.dataa(!\del_np_cnt[1]~q ),
	.datab(!\del_np_cnt[0]~q ),
	.datac(!\del_np_cnt[2]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_np_cnt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_np_cnt~5 .extended_lut = "off";
defparam \del_np_cnt~5 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \del_np_cnt~5 .shared_arith = "off";

dffeas \del_np_cnt[1] (
	.clk(clk),
	.d(\del_np_cnt~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_np_cnt[1]~q ),
	.prn(vcc));
defparam \del_np_cnt[1] .is_wysiwyg = "true";
defparam \del_np_cnt[1] .power_up = "low";

cyclonev_lcell_comb \del_np_cnt~4 (
	.dataa(!\del_np_cnt[2]~q ),
	.datab(!\del_np_cnt[1]~q ),
	.datac(!\del_np_cnt[0]~q ),
	.datad(!\del_np_cnt[2]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_np_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_np_cnt~4 .extended_lut = "off";
defparam \del_np_cnt~4 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \del_np_cnt~4 .shared_arith = "off";

dffeas \del_np_cnt[2] (
	.clk(clk),
	.d(\del_np_cnt~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_np_cnt[2]~q ),
	.prn(vcc));
defparam \del_np_cnt[2] .is_wysiwyg = "true";
defparam \del_np_cnt[2] .power_up = "low";

cyclonev_lcell_comb \del_np_cnt~3 (
	.dataa(!\del_np_cnt[3]~q ),
	.datab(!\del_np_cnt[2]~q ),
	.datac(!\del_np_cnt[1]~q ),
	.datad(!\del_np_cnt[0]~q ),
	.datae(!\del_np_cnt[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_np_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_np_cnt~3 .extended_lut = "off";
defparam \del_np_cnt~3 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \del_np_cnt~3 .shared_arith = "off";

dffeas \del_np_cnt[3] (
	.clk(clk),
	.d(\del_np_cnt~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_np_cnt[3]~q ),
	.prn(vcc));
defparam \del_np_cnt[3] .is_wysiwyg = "true";
defparam \del_np_cnt[3] .power_up = "low";

cyclonev_lcell_comb \del_np_cnt~2 (
	.dataa(!\del_np_cnt[4]~q ),
	.datab(!\del_np_cnt[3]~q ),
	.datac(!\del_np_cnt[2]~q ),
	.datad(!\del_np_cnt[1]~q ),
	.datae(!\del_np_cnt[0]~q ),
	.dataf(!\del_np_cnt[2]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_np_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_np_cnt~2 .extended_lut = "off";
defparam \del_np_cnt~2 .lut_mask = 64'h96696996FFFFFFFF;
defparam \del_np_cnt~2 .shared_arith = "off";

dffeas \del_np_cnt[4] (
	.clk(clk),
	.d(\del_np_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_np_cnt[4]~q ),
	.prn(vcc));
defparam \del_np_cnt[4] .is_wysiwyg = "true";
defparam \del_np_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\del_np_cnt[4]~q ),
	.datab(!\del_np_cnt[3]~q ),
	.datac(!\del_np_cnt[2]~q ),
	.datad(!\del_np_cnt[1]~q ),
	.datae(!\del_np_cnt[0]~q ),
	.dataf(!\sdetd.DISABLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!\sdetd.BLOCK_READY~q ),
	.datab(!\del_np_cnt[4]~q ),
	.datac(!\del_np_cnt[3]~q ),
	.datad(!\del_np_cnt[2]~q ),
	.datae(!\del_np_cnt[1]~q ),
	.dataf(!\del_np_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!\sdetd.ENABLE~q ),
	.datab(!\gen_blk_float:gen_streaming:gen_disc:delay_next_blk|tdl_arr[0]~q ),
	.datac(!\gen_blk_float:gen_streaming:gen_disc:gen_consts_64:delay_next_pass|tdl_arr[6]~q ),
	.datad(!\sdetd.IDLE~q ),
	.datae(!\Selector1~0_combout ),
	.dataf(!\Selector1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \Selector1~2 .shared_arith = "off";

dffeas \sdetd.ENABLE (
	.clk(clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sdetd.ENABLE~q ),
	.prn(vcc));
defparam \sdetd.ENABLE .is_wysiwyg = "true";
defparam \sdetd.ENABLE .power_up = "low";

cyclonev_lcell_comb \sdetd~8 (
	.dataa(!reset_n),
	.datab(!\sdetd.ENABLE~q ),
	.datac(!\gen_blk_float:gen_streaming:gen_disc:gen_consts_64:delay_next_pass|tdl_arr[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdetd~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdetd~8 .extended_lut = "off";
defparam \sdetd~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \sdetd~8 .shared_arith = "off";

dffeas \sdetd.GBLK (
	.clk(clk),
	.d(\sdetd~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sdetd.GBLK~q ),
	.prn(vcc));
defparam \sdetd.GBLK .is_wysiwyg = "true";
defparam \sdetd.GBLK .power_up = "low";

cyclonev_lcell_comb \gain_lut_8pts~0 (
	.dataa(!tdl_arr_3_1),
	.datab(!tdl_arr_7_1),
	.datac(!tdl_arr_3_11),
	.datad(!tdl_arr_7_11),
	.datae(!tdl_arr_3_12),
	.dataf(!tdl_arr_7_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~0 .extended_lut = "off";
defparam \gain_lut_8pts~0 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~0 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~1 (
	.dataa(!reg_no_twiddle603),
	.datab(!reg_no_twiddle607),
	.datac(!reg_no_twiddle617),
	.datad(!reg_no_twiddle613),
	.datae(!tdl_arr_3_13),
	.dataf(!tdl_arr_7_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~1 .extended_lut = "off";
defparam \gain_lut_8pts~1 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~1 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~2 (
	.dataa(!tdl_arr_3_14),
	.datab(!tdl_arr_7_14),
	.datac(!tdl_arr_3_15),
	.datad(!tdl_arr_7_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~2 .extended_lut = "off";
defparam \gain_lut_8pts~2 .lut_mask = 64'h6996699669966996;
defparam \gain_lut_8pts~2 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~3 (
	.dataa(!\sdetd.GBLK~q ),
	.datab(!\sdetd.ENABLE~q ),
	.datac(!\gain_lut_8pts~0_combout ),
	.datad(!\gain_lut_8pts~1_combout ),
	.datae(!\gain_lut_8pts~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~3 .extended_lut = "off";
defparam \gain_lut_8pts~3 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \gain_lut_8pts~3 .shared_arith = "off";

dffeas \gain_lut_8pts[0] (
	.clk(clk),
	.d(\gain_lut_8pts~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_8pts[0]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[0] .is_wysiwyg = "true";
defparam \gain_lut_8pts[0] .power_up = "low";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!\gain_lut_8pts[0]~q ),
	.datab(!\gain_lut_blk[0]~q ),
	.datac(!\sdetd.GBLK~q ),
	.datad(!\sdetd.ENABLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector6~0 .shared_arith = "off";

dffeas \gain_lut_blk[0] (
	.clk(clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_blk[0]~q ),
	.prn(vcc));
defparam \gain_lut_blk[0] .is_wysiwyg = "true";
defparam \gain_lut_blk[0] .power_up = "low";

cyclonev_lcell_comb \slb_i[0] (
	.dataa(!\gain_lut_8pts[0]~q ),
	.datab(!\gain_lut_blk[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_i[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_i[0] .extended_lut = "off";
defparam \slb_i[0] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \slb_i[0] .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~4 (
	.dataa(!tdl_arr_7_1),
	.datab(!tdl_arr_7_11),
	.datac(!tdl_arr_7_12),
	.datad(!tdl_arr_4_1),
	.datae(!tdl_arr_4_11),
	.dataf(!tdl_arr_4_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~4 .extended_lut = "off";
defparam \gain_lut_8pts~4 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~4 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~5 (
	.dataa(!reg_no_twiddle607),
	.datab(!reg_no_twiddle617),
	.datac(!tdl_arr_7_13),
	.datad(!reg_no_twiddle604),
	.datae(!reg_no_twiddle614),
	.dataf(!tdl_arr_4_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~5 .extended_lut = "off";
defparam \gain_lut_8pts~5 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~5 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~6 (
	.dataa(!tdl_arr_7_14),
	.datab(!tdl_arr_7_15),
	.datac(!tdl_arr_4_14),
	.datad(!tdl_arr_4_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~6 .extended_lut = "off";
defparam \gain_lut_8pts~6 .lut_mask = 64'h6996699669966996;
defparam \gain_lut_8pts~6 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~7 (
	.dataa(!\sdetd.GBLK~q ),
	.datab(!\sdetd.ENABLE~q ),
	.datac(!\gain_lut_8pts~4_combout ),
	.datad(!\gain_lut_8pts~5_combout ),
	.datae(!\gain_lut_8pts~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~7 .extended_lut = "off";
defparam \gain_lut_8pts~7 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \gain_lut_8pts~7 .shared_arith = "off";

dffeas \gain_lut_8pts[1] (
	.clk(clk),
	.d(\gain_lut_8pts~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_8pts[1]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[1] .is_wysiwyg = "true";
defparam \gain_lut_8pts[1] .power_up = "low";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!\gain_lut_8pts[1]~q ),
	.datab(!\gain_lut_blk[1]~q ),
	.datac(!\sdetd.GBLK~q ),
	.datad(!\sdetd.ENABLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector5~0 .shared_arith = "off";

dffeas \gain_lut_blk[1] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_blk[1]~q ),
	.prn(vcc));
defparam \gain_lut_blk[1] .is_wysiwyg = "true";
defparam \gain_lut_blk[1] .power_up = "low";

cyclonev_lcell_comb \slb_i[1] (
	.dataa(!\gain_lut_8pts[1]~q ),
	.datab(!\gain_lut_blk[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_i[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_i[1] .extended_lut = "off";
defparam \slb_i[1] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \slb_i[1] .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~8 (
	.dataa(!tdl_arr_7_1),
	.datab(!tdl_arr_7_11),
	.datac(!tdl_arr_7_12),
	.datad(!tdl_arr_5_1),
	.datae(!tdl_arr_5_11),
	.dataf(!tdl_arr_5_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~8 .extended_lut = "off";
defparam \gain_lut_8pts~8 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~8 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~9 (
	.dataa(!reg_no_twiddle607),
	.datab(!reg_no_twiddle617),
	.datac(!tdl_arr_7_13),
	.datad(!reg_no_twiddle605),
	.datae(!reg_no_twiddle615),
	.dataf(!tdl_arr_5_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~9 .extended_lut = "off";
defparam \gain_lut_8pts~9 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~9 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~10 (
	.dataa(!tdl_arr_7_14),
	.datab(!tdl_arr_7_15),
	.datac(!tdl_arr_5_14),
	.datad(!tdl_arr_5_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~10 .extended_lut = "off";
defparam \gain_lut_8pts~10 .lut_mask = 64'h6996699669966996;
defparam \gain_lut_8pts~10 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~11 (
	.dataa(!\sdetd.GBLK~q ),
	.datab(!\sdetd.ENABLE~q ),
	.datac(!\gain_lut_8pts~8_combout ),
	.datad(!\gain_lut_8pts~9_combout ),
	.datae(!\gain_lut_8pts~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~11 .extended_lut = "off";
defparam \gain_lut_8pts~11 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \gain_lut_8pts~11 .shared_arith = "off";

dffeas \gain_lut_8pts[2] (
	.clk(clk),
	.d(\gain_lut_8pts~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_8pts[2]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[2] .is_wysiwyg = "true";
defparam \gain_lut_8pts[2] .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!\gain_lut_8pts[2]~q ),
	.datab(!\gain_lut_blk[2]~q ),
	.datac(!\sdetd.GBLK~q ),
	.datad(!\sdetd.ENABLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector4~0 .shared_arith = "off";

dffeas \gain_lut_blk[2] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_blk[2]~q ),
	.prn(vcc));
defparam \gain_lut_blk[2] .is_wysiwyg = "true";
defparam \gain_lut_blk[2] .power_up = "low";

cyclonev_lcell_comb \slb_i[2] (
	.dataa(!\gain_lut_8pts[2]~q ),
	.datab(!\gain_lut_blk[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_i[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_i[2] .extended_lut = "off";
defparam \slb_i[2] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \slb_i[2] .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~12 (
	.dataa(!tdl_arr_7_1),
	.datab(!tdl_arr_7_11),
	.datac(!tdl_arr_7_12),
	.datad(!tdl_arr_6_1),
	.datae(!tdl_arr_6_11),
	.dataf(!tdl_arr_6_12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~12 .extended_lut = "off";
defparam \gain_lut_8pts~12 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~12 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~13 (
	.dataa(!reg_no_twiddle607),
	.datab(!reg_no_twiddle617),
	.datac(!tdl_arr_7_13),
	.datad(!reg_no_twiddle606),
	.datae(!reg_no_twiddle616),
	.dataf(!tdl_arr_6_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~13 .extended_lut = "off";
defparam \gain_lut_8pts~13 .lut_mask = 64'h6996966996696996;
defparam \gain_lut_8pts~13 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~14 (
	.dataa(!tdl_arr_7_14),
	.datab(!tdl_arr_7_15),
	.datac(!tdl_arr_6_14),
	.datad(!tdl_arr_6_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~14 .extended_lut = "off";
defparam \gain_lut_8pts~14 .lut_mask = 64'h6996699669966996;
defparam \gain_lut_8pts~14 .shared_arith = "off";

cyclonev_lcell_comb \gain_lut_8pts~15 (
	.dataa(!\sdetd.GBLK~q ),
	.datab(!\sdetd.ENABLE~q ),
	.datac(!\gain_lut_8pts~12_combout ),
	.datad(!\gain_lut_8pts~13_combout ),
	.datae(!\gain_lut_8pts~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gain_lut_8pts~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gain_lut_8pts~15 .extended_lut = "off";
defparam \gain_lut_8pts~15 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \gain_lut_8pts~15 .shared_arith = "off";

dffeas \gain_lut_8pts[3] (
	.clk(clk),
	.d(\gain_lut_8pts~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_8pts[3]~q ),
	.prn(vcc));
defparam \gain_lut_8pts[3] .is_wysiwyg = "true";
defparam \gain_lut_8pts[3] .power_up = "low";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\gain_lut_8pts[3]~q ),
	.datab(!\gain_lut_blk[3]~q ),
	.datac(!\sdetd.GBLK~q ),
	.datad(!\sdetd.ENABLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector3~0 .shared_arith = "off";

dffeas \gain_lut_blk[3] (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\gain_lut_blk[3]~q ),
	.prn(vcc));
defparam \gain_lut_blk[3] .is_wysiwyg = "true";
defparam \gain_lut_blk[3] .power_up = "low";

cyclonev_lcell_comb \slb_i[3] (
	.dataa(!\gain_lut_8pts[3]~q ),
	.datab(!\gain_lut_blk[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\slb_i[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \slb_i[3] .extended_lut = "off";
defparam \slb_i[3] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \slb_i[3] .shared_arith = "off";

cyclonev_lcell_comb \lut_out_tmp~0 (
	.dataa(!\slb_i[0]~combout ),
	.datab(!\slb_i[1]~combout ),
	.datac(!\slb_i[2]~combout ),
	.datad(!\slb_i[3]~combout ),
	.datae(!reset_n),
	.dataf(!\sdetd.SLBI~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lut_out_tmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lut_out_tmp~0 .extended_lut = "off";
defparam \lut_out_tmp~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \lut_out_tmp~0 .shared_arith = "off";

cyclonev_lcell_comb \lut_out_tmp[2]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\sdetd.SLBI~q ),
	.datad(!\sdetd.BLOCK_READY~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lut_out_tmp[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lut_out_tmp[2]~1 .extended_lut = "off";
defparam \lut_out_tmp[2]~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \lut_out_tmp[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \lut_out_tmp~2 (
	.dataa(!\slb_i[0]~combout ),
	.datab(!\slb_i[1]~combout ),
	.datac(!\slb_i[2]~combout ),
	.datad(!\slb_i[3]~combout ),
	.datae(!reset_n),
	.dataf(!\sdetd.SLBI~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lut_out_tmp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lut_out_tmp~2 .extended_lut = "off";
defparam \lut_out_tmp~2 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \lut_out_tmp~2 .shared_arith = "off";

cyclonev_lcell_comb \lut_out_tmp~3 (
	.dataa(!reset_n),
	.datab(!\slb_i[0]~combout ),
	.datac(!\slb_i[1]~combout ),
	.datad(!\slb_i[2]~combout ),
	.datae(!\slb_i[3]~combout ),
	.dataf(!\sdetd.SLBI~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lut_out_tmp~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lut_out_tmp~3 .extended_lut = "off";
defparam \lut_out_tmp~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \lut_out_tmp~3 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl_bit_rst_2 (
	next_block,
	tdl_arr_0,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	next_block;
output 	tdl_arr_0;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \tdl_arr[0] (
	.clk(clk),
	.d(next_block),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_bit_rst_3 (
	tdl_arr_6,
	tdl_arr_9,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_6;
input 	tdl_arr_9;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;


dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_6),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(tdl_arr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

endmodule

module IFFT_asj_fft_pround_6 (
	butterfly_st2006,
	butterfly_st2009,
	butterfly_st2007,
	butterfly_st2008,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	global_clock_enable,
	pipeline_dffe_6,
	pipeline_dffe_9,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2006;
input 	butterfly_st2009;
input 	butterfly_st2007;
input 	butterfly_st2008;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	global_clock_enable;
output 	pipeline_dffe_6;
output 	pipeline_dffe_9;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_7 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2006(butterfly_st2006),
	.butterfly_st2009(butterfly_st2009),
	.butterfly_st2007(butterfly_st2007),
	.butterfly_st2008(butterfly_st2008),
	.butterfly_st2005(butterfly_st2005),
	.butterfly_st2004(butterfly_st2004),
	.butterfly_st2003(butterfly_st2003),
	.butterfly_st2002(butterfly_st2002),
	.butterfly_st2001(butterfly_st2001),
	.butterfly_st2000(butterfly_st2000),
	.clken(global_clock_enable),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_7 (
	butterfly_st2006,
	butterfly_st2009,
	butterfly_st2007,
	butterfly_st2008,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	clken,
	pipeline_dffe_6,
	pipeline_dffe_9,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2006;
input 	butterfly_st2009;
input 	butterfly_st2007;
input 	butterfly_st2008;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	clken;
output 	pipeline_dffe_6;
output 	pipeline_dffe_9;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj auto_generated(
	.butterfly_st2006(butterfly_st2006),
	.butterfly_st2009(butterfly_st2009),
	.butterfly_st2007(butterfly_st2007),
	.butterfly_st2008(butterfly_st2008),
	.butterfly_st2005(butterfly_st2005),
	.butterfly_st2004(butterfly_st2004),
	.butterfly_st2003(butterfly_st2003),
	.butterfly_st2002(butterfly_st2002),
	.butterfly_st2001(butterfly_st2001),
	.butterfly_st2000(butterfly_st2000),
	.clken(clken),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj (
	butterfly_st2006,
	butterfly_st2009,
	butterfly_st2007,
	butterfly_st2008,
	butterfly_st2005,
	butterfly_st2004,
	butterfly_st2003,
	butterfly_st2002,
	butterfly_st2001,
	butterfly_st2000,
	clken,
	pipeline_dffe_6,
	pipeline_dffe_9,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2006;
input 	butterfly_st2009;
input 	butterfly_st2007;
input 	butterfly_st2008;
input 	butterfly_st2005;
input 	butterfly_st2004;
input 	butterfly_st2003;
input 	butterfly_st2002;
input 	butterfly_st2001;
input 	butterfly_st2000;
input 	clken;
output 	pipeline_dffe_6;
output 	pipeline_dffe_9;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2009),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2000),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2001),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2002),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2003),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2004),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2005),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2006),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2007),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2008),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2009),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_7 (
	butterfly_st2019,
	butterfly_st2016,
	butterfly_st2017,
	butterfly_st2018,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	global_clock_enable,
	pipeline_dffe_9,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2019;
input 	butterfly_st2016;
input 	butterfly_st2017;
input 	butterfly_st2018;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	global_clock_enable;
output 	pipeline_dffe_9;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_8 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2019(butterfly_st2019),
	.butterfly_st2016(butterfly_st2016),
	.butterfly_st2017(butterfly_st2017),
	.butterfly_st2018(butterfly_st2018),
	.butterfly_st2015(butterfly_st2015),
	.butterfly_st2014(butterfly_st2014),
	.butterfly_st2013(butterfly_st2013),
	.butterfly_st2012(butterfly_st2012),
	.butterfly_st2011(butterfly_st2011),
	.butterfly_st2010(butterfly_st2010),
	.clken(global_clock_enable),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_8 (
	butterfly_st2019,
	butterfly_st2016,
	butterfly_st2017,
	butterfly_st2018,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	clken,
	pipeline_dffe_9,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2019;
input 	butterfly_st2016;
input 	butterfly_st2017;
input 	butterfly_st2018;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	clken;
output 	pipeline_dffe_9;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_1 auto_generated(
	.butterfly_st2019(butterfly_st2019),
	.butterfly_st2016(butterfly_st2016),
	.butterfly_st2017(butterfly_st2017),
	.butterfly_st2018(butterfly_st2018),
	.butterfly_st2015(butterfly_st2015),
	.butterfly_st2014(butterfly_st2014),
	.butterfly_st2013(butterfly_st2013),
	.butterfly_st2012(butterfly_st2012),
	.butterfly_st2011(butterfly_st2011),
	.butterfly_st2010(butterfly_st2010),
	.clken(clken),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_1 (
	butterfly_st2019,
	butterfly_st2016,
	butterfly_st2017,
	butterfly_st2018,
	butterfly_st2015,
	butterfly_st2014,
	butterfly_st2013,
	butterfly_st2012,
	butterfly_st2011,
	butterfly_st2010,
	clken,
	pipeline_dffe_9,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2019;
input 	butterfly_st2016;
input 	butterfly_st2017;
input 	butterfly_st2018;
input 	butterfly_st2015;
input 	butterfly_st2014;
input 	butterfly_st2013;
input 	butterfly_st2012;
input 	butterfly_st2011;
input 	butterfly_st2010;
input 	clken;
output 	pipeline_dffe_9;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2019),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2010),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2011),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2012),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2013),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2014),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2015),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2016),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2017),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2018),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2019),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:0:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_8 (
	butterfly_st2102,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	butterfly_st2109,
	butterfly_st2101,
	butterfly_st2100,
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2102;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	butterfly_st2109;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_9 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2102(butterfly_st2102),
	.butterfly_st2103(butterfly_st2103),
	.butterfly_st2104(butterfly_st2104),
	.butterfly_st2105(butterfly_st2105),
	.butterfly_st2106(butterfly_st2106),
	.butterfly_st2107(butterfly_st2107),
	.butterfly_st2108(butterfly_st2108),
	.butterfly_st2109(butterfly_st2109),
	.butterfly_st2101(butterfly_st2101),
	.butterfly_st2100(butterfly_st2100),
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_9 (
	butterfly_st2102,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	butterfly_st2109,
	butterfly_st2101,
	butterfly_st2100,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2102;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	butterfly_st2109;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_2 auto_generated(
	.butterfly_st2102(butterfly_st2102),
	.butterfly_st2103(butterfly_st2103),
	.butterfly_st2104(butterfly_st2104),
	.butterfly_st2105(butterfly_st2105),
	.butterfly_st2106(butterfly_st2106),
	.butterfly_st2107(butterfly_st2107),
	.butterfly_st2108(butterfly_st2108),
	.butterfly_st2109(butterfly_st2109),
	.butterfly_st2101(butterfly_st2101),
	.butterfly_st2100(butterfly_st2100),
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_2 (
	butterfly_st2102,
	butterfly_st2103,
	butterfly_st2104,
	butterfly_st2105,
	butterfly_st2106,
	butterfly_st2107,
	butterfly_st2108,
	butterfly_st2109,
	butterfly_st2101,
	butterfly_st2100,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2102;
input 	butterfly_st2103;
input 	butterfly_st2104;
input 	butterfly_st2105;
input 	butterfly_st2106;
input 	butterfly_st2107;
input 	butterfly_st2108;
input 	butterfly_st2109;
input 	butterfly_st2101;
input 	butterfly_st2100;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2109),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2100),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2102),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2103),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2104),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2105),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2106),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2107),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2108),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2109),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_9 (
	butterfly_st2112,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	butterfly_st2119,
	butterfly_st2111,
	butterfly_st2110,
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2112;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	butterfly_st2119;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_10 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2112(butterfly_st2112),
	.butterfly_st2113(butterfly_st2113),
	.butterfly_st2114(butterfly_st2114),
	.butterfly_st2115(butterfly_st2115),
	.butterfly_st2116(butterfly_st2116),
	.butterfly_st2117(butterfly_st2117),
	.butterfly_st2118(butterfly_st2118),
	.butterfly_st2119(butterfly_st2119),
	.butterfly_st2111(butterfly_st2111),
	.butterfly_st2110(butterfly_st2110),
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_10 (
	butterfly_st2112,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	butterfly_st2119,
	butterfly_st2111,
	butterfly_st2110,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2112;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	butterfly_st2119;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_3 auto_generated(
	.butterfly_st2112(butterfly_st2112),
	.butterfly_st2113(butterfly_st2113),
	.butterfly_st2114(butterfly_st2114),
	.butterfly_st2115(butterfly_st2115),
	.butterfly_st2116(butterfly_st2116),
	.butterfly_st2117(butterfly_st2117),
	.butterfly_st2118(butterfly_st2118),
	.butterfly_st2119(butterfly_st2119),
	.butterfly_st2111(butterfly_st2111),
	.butterfly_st2110(butterfly_st2110),
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_3 (
	butterfly_st2112,
	butterfly_st2113,
	butterfly_st2114,
	butterfly_st2115,
	butterfly_st2116,
	butterfly_st2117,
	butterfly_st2118,
	butterfly_st2119,
	butterfly_st2111,
	butterfly_st2110,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2112;
input 	butterfly_st2113;
input 	butterfly_st2114;
input 	butterfly_st2115;
input 	butterfly_st2116;
input 	butterfly_st2117;
input 	butterfly_st2118;
input 	butterfly_st2119;
input 	butterfly_st2111;
input 	butterfly_st2110;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2119),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2112),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2113),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2114),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2115),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2116),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2117),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2118),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2119),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:1:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_10 (
	butterfly_st2202,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	butterfly_st2209,
	butterfly_st2201,
	butterfly_st2200,
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2202;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	butterfly_st2209;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_11 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2202(butterfly_st2202),
	.butterfly_st2203(butterfly_st2203),
	.butterfly_st2204(butterfly_st2204),
	.butterfly_st2205(butterfly_st2205),
	.butterfly_st2206(butterfly_st2206),
	.butterfly_st2207(butterfly_st2207),
	.butterfly_st2208(butterfly_st2208),
	.butterfly_st2209(butterfly_st2209),
	.butterfly_st2201(butterfly_st2201),
	.butterfly_st2200(butterfly_st2200),
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_11 (
	butterfly_st2202,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	butterfly_st2209,
	butterfly_st2201,
	butterfly_st2200,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2202;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	butterfly_st2209;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_4 auto_generated(
	.butterfly_st2202(butterfly_st2202),
	.butterfly_st2203(butterfly_st2203),
	.butterfly_st2204(butterfly_st2204),
	.butterfly_st2205(butterfly_st2205),
	.butterfly_st2206(butterfly_st2206),
	.butterfly_st2207(butterfly_st2207),
	.butterfly_st2208(butterfly_st2208),
	.butterfly_st2209(butterfly_st2209),
	.butterfly_st2201(butterfly_st2201),
	.butterfly_st2200(butterfly_st2200),
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_4 (
	butterfly_st2202,
	butterfly_st2203,
	butterfly_st2204,
	butterfly_st2205,
	butterfly_st2206,
	butterfly_st2207,
	butterfly_st2208,
	butterfly_st2209,
	butterfly_st2201,
	butterfly_st2200,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2202;
input 	butterfly_st2203;
input 	butterfly_st2204;
input 	butterfly_st2205;
input 	butterfly_st2206;
input 	butterfly_st2207;
input 	butterfly_st2208;
input 	butterfly_st2209;
input 	butterfly_st2201;
input 	butterfly_st2200;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2209),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2200),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2201),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2202),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2203),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2204),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2205),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2206),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2207),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2208),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2209),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_11 (
	butterfly_st2212,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	butterfly_st2219,
	butterfly_st2211,
	butterfly_st2210,
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2212;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	butterfly_st2219;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_12 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2212(butterfly_st2212),
	.butterfly_st2213(butterfly_st2213),
	.butterfly_st2214(butterfly_st2214),
	.butterfly_st2215(butterfly_st2215),
	.butterfly_st2216(butterfly_st2216),
	.butterfly_st2217(butterfly_st2217),
	.butterfly_st2218(butterfly_st2218),
	.butterfly_st2219(butterfly_st2219),
	.butterfly_st2211(butterfly_st2211),
	.butterfly_st2210(butterfly_st2210),
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_12 (
	butterfly_st2212,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	butterfly_st2219,
	butterfly_st2211,
	butterfly_st2210,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2212;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	butterfly_st2219;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_5 auto_generated(
	.butterfly_st2212(butterfly_st2212),
	.butterfly_st2213(butterfly_st2213),
	.butterfly_st2214(butterfly_st2214),
	.butterfly_st2215(butterfly_st2215),
	.butterfly_st2216(butterfly_st2216),
	.butterfly_st2217(butterfly_st2217),
	.butterfly_st2218(butterfly_st2218),
	.butterfly_st2219(butterfly_st2219),
	.butterfly_st2211(butterfly_st2211),
	.butterfly_st2210(butterfly_st2210),
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_5 (
	butterfly_st2212,
	butterfly_st2213,
	butterfly_st2214,
	butterfly_st2215,
	butterfly_st2216,
	butterfly_st2217,
	butterfly_st2218,
	butterfly_st2219,
	butterfly_st2211,
	butterfly_st2210,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2212;
input 	butterfly_st2213;
input 	butterfly_st2214;
input 	butterfly_st2215;
input 	butterfly_st2216;
input 	butterfly_st2217;
input 	butterfly_st2218;
input 	butterfly_st2219;
input 	butterfly_st2211;
input 	butterfly_st2210;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2219),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2210),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2211),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2212),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2213),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2214),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2215),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2216),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2217),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2218),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2219),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:2:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_12 (
	butterfly_st2302,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	butterfly_st2309,
	butterfly_st2301,
	butterfly_st2300,
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2302;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	butterfly_st2309;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_13 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2302(butterfly_st2302),
	.butterfly_st2303(butterfly_st2303),
	.butterfly_st2304(butterfly_st2304),
	.butterfly_st2305(butterfly_st2305),
	.butterfly_st2306(butterfly_st2306),
	.butterfly_st2307(butterfly_st2307),
	.butterfly_st2308(butterfly_st2308),
	.butterfly_st2309(butterfly_st2309),
	.butterfly_st2301(butterfly_st2301),
	.butterfly_st2300(butterfly_st2300),
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_13 (
	butterfly_st2302,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	butterfly_st2309,
	butterfly_st2301,
	butterfly_st2300,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2302;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	butterfly_st2309;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_6 auto_generated(
	.butterfly_st2302(butterfly_st2302),
	.butterfly_st2303(butterfly_st2303),
	.butterfly_st2304(butterfly_st2304),
	.butterfly_st2305(butterfly_st2305),
	.butterfly_st2306(butterfly_st2306),
	.butterfly_st2307(butterfly_st2307),
	.butterfly_st2308(butterfly_st2308),
	.butterfly_st2309(butterfly_st2309),
	.butterfly_st2301(butterfly_st2301),
	.butterfly_st2300(butterfly_st2300),
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_6 (
	butterfly_st2302,
	butterfly_st2303,
	butterfly_st2304,
	butterfly_st2305,
	butterfly_st2306,
	butterfly_st2307,
	butterfly_st2308,
	butterfly_st2309,
	butterfly_st2301,
	butterfly_st2300,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2302;
input 	butterfly_st2303;
input 	butterfly_st2304;
input 	butterfly_st2305;
input 	butterfly_st2306;
input 	butterfly_st2307;
input 	butterfly_st2308;
input 	butterfly_st2309;
input 	butterfly_st2301;
input 	butterfly_st2300;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2309),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2300),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2301),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2302),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2303),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2304),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2305),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2306),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2307),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2308),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2309),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_13 (
	butterfly_st2312,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	butterfly_st2319,
	butterfly_st2311,
	butterfly_st2310,
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2312;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	butterfly_st2319;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_14 \gbrnd:nev:gp:lpm_add_sub_component (
	.butterfly_st2312(butterfly_st2312),
	.butterfly_st2313(butterfly_st2313),
	.butterfly_st2314(butterfly_st2314),
	.butterfly_st2315(butterfly_st2315),
	.butterfly_st2316(butterfly_st2316),
	.butterfly_st2317(butterfly_st2317),
	.butterfly_st2318(butterfly_st2318),
	.butterfly_st2319(butterfly_st2319),
	.butterfly_st2311(butterfly_st2311),
	.butterfly_st2310(butterfly_st2310),
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_14 (
	butterfly_st2312,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	butterfly_st2319,
	butterfly_st2311,
	butterfly_st2310,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2312;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	butterfly_st2319;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_7 auto_generated(
	.butterfly_st2312(butterfly_st2312),
	.butterfly_st2313(butterfly_st2313),
	.butterfly_st2314(butterfly_st2314),
	.butterfly_st2315(butterfly_st2315),
	.butterfly_st2316(butterfly_st2316),
	.butterfly_st2317(butterfly_st2317),
	.butterfly_st2318(butterfly_st2318),
	.butterfly_st2319(butterfly_st2319),
	.butterfly_st2311(butterfly_st2311),
	.butterfly_st2310(butterfly_st2310),
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_7 (
	butterfly_st2312,
	butterfly_st2313,
	butterfly_st2314,
	butterfly_st2315,
	butterfly_st2316,
	butterfly_st2317,
	butterfly_st2318,
	butterfly_st2319,
	butterfly_st2311,
	butterfly_st2310,
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock)/* synthesis synthesis_greybox=1 */;
input 	butterfly_st2312;
input 	butterfly_st2313;
input 	butterfly_st2314;
input 	butterfly_st2315;
input 	butterfly_st2316;
input 	butterfly_st2317;
input 	butterfly_st2318;
input 	butterfly_st2319;
input 	butterfly_st2311;
input 	butterfly_st2310;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2319),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2310),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2311),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2312),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2313),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2314),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2315),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2316),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2317),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2318),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!butterfly_st2319),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_dft_1:bfpdft|gen_full_rnd:gen_rounding_blk:3:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_in_write_sgl (
	next_block1,
	data_rdy_int1,
	wren_1,
	data_in_r_6,
	wr_address_i_int_0,
	wr_address_i_int_1,
	wr_address_i_int_2,
	wr_address_i_int_3,
	wren_2,
	wren_3,
	wren_0,
	data_in_r_5,
	data_in_r_2,
	data_in_r_3,
	data_in_r_4,
	data_in_r_7,
	data_in_i_7,
	data_in_i_6,
	data_in_i_3,
	data_in_i_4,
	data_in_i_5,
	data_in_i_2,
	data_in_r_0,
	data_in_r_1,
	data_in_i_0,
	data_in_i_1,
	core_real_in_6,
	core_real_in_5,
	core_real_in_2,
	core_real_in_3,
	core_real_in_4,
	core_real_in_7,
	core_imag_in_7,
	core_imag_in_6,
	core_imag_in_3,
	core_imag_in_4,
	core_imag_in_5,
	core_imag_in_2,
	core_real_in_0,
	core_real_in_1,
	core_imag_in_0,
	core_imag_in_1,
	anb1,
	send_sop_s,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	next_block1;
output 	data_rdy_int1;
output 	wren_1;
output 	data_in_r_6;
output 	wr_address_i_int_0;
output 	wr_address_i_int_1;
output 	wr_address_i_int_2;
output 	wr_address_i_int_3;
output 	wren_2;
output 	wren_3;
output 	wren_0;
output 	data_in_r_5;
output 	data_in_r_2;
output 	data_in_r_3;
output 	data_in_r_4;
output 	data_in_r_7;
output 	data_in_i_7;
output 	data_in_i_6;
output 	data_in_i_3;
output 	data_in_i_4;
output 	data_in_i_5;
output 	data_in_i_2;
output 	data_in_r_0;
output 	data_in_r_1;
output 	data_in_i_0;
output 	data_in_i_1;
input 	core_real_in_6;
input 	core_real_in_5;
input 	core_real_in_2;
input 	core_real_in_3;
input 	core_real_in_4;
input 	core_real_in_7;
input 	core_imag_in_7;
input 	core_imag_in_6;
input 	core_imag_in_3;
input 	core_imag_in_4;
input 	core_imag_in_5;
input 	core_imag_in_2;
input 	core_real_in_0;
input 	core_real_in_1;
input 	core_imag_in_0;
input 	core_imag_in_1;
output 	anb1;
input 	send_sop_s;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \str_count_en~0_combout ;
wire \str_count_en~q ;
wire \Add0~17_sumout ;
wire \counter_i~0_combout ;
wire \count[0]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \count[1]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \count[2]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \count[3]~q ;
wire \Add0~10 ;
wire \Add0~21_sumout ;
wire \count[4]~q ;
wire \Add0~22 ;
wire \Add0~13_sumout ;
wire \count[5]~q ;
wire \Equal0~0_combout ;
wire \data_rdy_int~0_combout ;
wire \Add1~0_combout ;
wire \sw[0]~q ;
wire \Add1~1_combout ;
wire \sw[1]~q ;
wire \Mux1~0_combout ;
wire \wr_addr[0]~q ;
wire \wr_addr[1]~q ;
wire \wr_addr[2]~q ;
wire \wr_addr[3]~q ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \Mux3~0_combout ;
wire \anb~0_combout ;


dffeas next_block(
	.clk(clk),
	.d(\Equal0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(next_block1),
	.prn(vcc));
defparam next_block.is_wysiwyg = "true";
defparam next_block.power_up = "low";

dffeas data_rdy_int(
	.clk(clk),
	.d(\data_rdy_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_rdy_int1),
	.prn(vcc));
defparam data_rdy_int.is_wysiwyg = "true";
defparam data_rdy_int.power_up = "low";

dffeas \wren[1] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wren_1),
	.prn(vcc));
defparam \wren[1] .is_wysiwyg = "true";
defparam \wren[1] .power_up = "low";

dffeas \data_in_r[6] (
	.clk(clk),
	.d(core_real_in_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_6),
	.prn(vcc));
defparam \data_in_r[6] .is_wysiwyg = "true";
defparam \data_in_r[6] .power_up = "low";

dffeas \wr_address_i_int[0] (
	.clk(clk),
	.d(\wr_addr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wr_address_i_int_0),
	.prn(vcc));
defparam \wr_address_i_int[0] .is_wysiwyg = "true";
defparam \wr_address_i_int[0] .power_up = "low";

dffeas \wr_address_i_int[1] (
	.clk(clk),
	.d(\wr_addr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wr_address_i_int_1),
	.prn(vcc));
defparam \wr_address_i_int[1] .is_wysiwyg = "true";
defparam \wr_address_i_int[1] .power_up = "low";

dffeas \wr_address_i_int[2] (
	.clk(clk),
	.d(\wr_addr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wr_address_i_int_2),
	.prn(vcc));
defparam \wr_address_i_int[2] .is_wysiwyg = "true";
defparam \wr_address_i_int[2] .power_up = "low";

dffeas \wr_address_i_int[3] (
	.clk(clk),
	.d(\wr_addr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wr_address_i_int_3),
	.prn(vcc));
defparam \wr_address_i_int[3] .is_wysiwyg = "true";
defparam \wr_address_i_int[3] .power_up = "low";

dffeas \wren[2] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wren_2),
	.prn(vcc));
defparam \wren[2] .is_wysiwyg = "true";
defparam \wren[2] .power_up = "low";

dffeas \wren[3] (
	.clk(clk),
	.d(\Mux1~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wren_3),
	.prn(vcc));
defparam \wren[3] .is_wysiwyg = "true";
defparam \wren[3] .power_up = "low";

dffeas \wren[0] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wren_0),
	.prn(vcc));
defparam \wren[0] .is_wysiwyg = "true";
defparam \wren[0] .power_up = "low";

dffeas \data_in_r[5] (
	.clk(clk),
	.d(core_real_in_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_5),
	.prn(vcc));
defparam \data_in_r[5] .is_wysiwyg = "true";
defparam \data_in_r[5] .power_up = "low";

dffeas \data_in_r[2] (
	.clk(clk),
	.d(core_real_in_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_2),
	.prn(vcc));
defparam \data_in_r[2] .is_wysiwyg = "true";
defparam \data_in_r[2] .power_up = "low";

dffeas \data_in_r[3] (
	.clk(clk),
	.d(core_real_in_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_3),
	.prn(vcc));
defparam \data_in_r[3] .is_wysiwyg = "true";
defparam \data_in_r[3] .power_up = "low";

dffeas \data_in_r[4] (
	.clk(clk),
	.d(core_real_in_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_4),
	.prn(vcc));
defparam \data_in_r[4] .is_wysiwyg = "true";
defparam \data_in_r[4] .power_up = "low";

dffeas \data_in_r[7] (
	.clk(clk),
	.d(core_real_in_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_7),
	.prn(vcc));
defparam \data_in_r[7] .is_wysiwyg = "true";
defparam \data_in_r[7] .power_up = "low";

dffeas \data_in_i[7] (
	.clk(clk),
	.d(core_imag_in_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_7),
	.prn(vcc));
defparam \data_in_i[7] .is_wysiwyg = "true";
defparam \data_in_i[7] .power_up = "low";

dffeas \data_in_i[6] (
	.clk(clk),
	.d(core_imag_in_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_6),
	.prn(vcc));
defparam \data_in_i[6] .is_wysiwyg = "true";
defparam \data_in_i[6] .power_up = "low";

dffeas \data_in_i[3] (
	.clk(clk),
	.d(core_imag_in_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_3),
	.prn(vcc));
defparam \data_in_i[3] .is_wysiwyg = "true";
defparam \data_in_i[3] .power_up = "low";

dffeas \data_in_i[4] (
	.clk(clk),
	.d(core_imag_in_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_4),
	.prn(vcc));
defparam \data_in_i[4] .is_wysiwyg = "true";
defparam \data_in_i[4] .power_up = "low";

dffeas \data_in_i[5] (
	.clk(clk),
	.d(core_imag_in_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_5),
	.prn(vcc));
defparam \data_in_i[5] .is_wysiwyg = "true";
defparam \data_in_i[5] .power_up = "low";

dffeas \data_in_i[2] (
	.clk(clk),
	.d(core_imag_in_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_2),
	.prn(vcc));
defparam \data_in_i[2] .is_wysiwyg = "true";
defparam \data_in_i[2] .power_up = "low";

dffeas \data_in_r[0] (
	.clk(clk),
	.d(core_real_in_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_0),
	.prn(vcc));
defparam \data_in_r[0] .is_wysiwyg = "true";
defparam \data_in_r[0] .power_up = "low";

dffeas \data_in_r[1] (
	.clk(clk),
	.d(core_real_in_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_r_1),
	.prn(vcc));
defparam \data_in_r[1] .is_wysiwyg = "true";
defparam \data_in_r[1] .power_up = "low";

dffeas \data_in_i[0] (
	.clk(clk),
	.d(core_imag_in_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_0),
	.prn(vcc));
defparam \data_in_i[0] .is_wysiwyg = "true";
defparam \data_in_i[0] .power_up = "low";

dffeas \data_in_i[1] (
	.clk(clk),
	.d(core_imag_in_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_in_i_1),
	.prn(vcc));
defparam \data_in_i[1] .is_wysiwyg = "true";
defparam \data_in_i[1] .power_up = "low";

dffeas anb(
	.clk(clk),
	.d(\anb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(!global_clock_enable),
	.q(anb1),
	.prn(vcc));
defparam anb.is_wysiwyg = "true";
defparam anb.power_up = "low";

cyclonev_lcell_comb \str_count_en~0 (
	.dataa(!send_sop_s),
	.datab(!\str_count_en~q ),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\str_count_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \str_count_en~0 .extended_lut = "off";
defparam \str_count_en~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \str_count_en~0 .shared_arith = "off";

dffeas str_count_en(
	.clk(clk),
	.d(\str_count_en~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\str_count_en~q ),
	.prn(vcc));
defparam str_count_en.is_wysiwyg = "true";
defparam str_count_en.power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\str_count_en~q ),
	.datae(gnd),
	.dataf(!\count[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \counter_i~0 (
	.dataa(!reset_n),
	.datab(!send_sop_s),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_i~0 .extended_lut = "off";
defparam \counter_i~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \counter_i~0 .shared_arith = "off";

dffeas \count[0] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \count[1] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \count[2] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \count[3] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \count[4] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \count[5] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\counter_i~0_combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\count[1]~q ),
	.datab(!\count[2]~q ),
	.datac(!\count[3]~q ),
	.datad(!\count[5]~q ),
	.datae(!\count[0]~q ),
	.dataf(!\count[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_rdy_int~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!data_rdy_int1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_rdy_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_rdy_int~0 .extended_lut = "off";
defparam \data_rdy_int~0 .lut_mask = 64'h7777777777777777;
defparam \data_rdy_int~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\count[0]~q ),
	.datab(!\count[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h6666666666666666;
defparam \Add1~0 .shared_arith = "off";

dffeas \sw[0] (
	.clk(clk),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw[0]~q ),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\count[1]~q ),
	.datab(!\count[5]~q ),
	.datac(!\count[0]~q ),
	.datad(!\count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6996699669966996;
defparam \Add1~1 .shared_arith = "off";

dffeas \sw[1] (
	.clk(clk),
	.d(\Add1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sw[1]~q ),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!\sw[0]~q ),
	.datab(!\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Mux1~0 .shared_arith = "off";

dffeas \wr_addr[0] (
	.clk(clk),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\wr_addr[0]~q ),
	.prn(vcc));
defparam \wr_addr[0] .is_wysiwyg = "true";
defparam \wr_addr[0] .power_up = "low";

dffeas \wr_addr[1] (
	.clk(clk),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\wr_addr[1]~q ),
	.prn(vcc));
defparam \wr_addr[1] .is_wysiwyg = "true";
defparam \wr_addr[1] .power_up = "low";

dffeas \wr_addr[2] (
	.clk(clk),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\wr_addr[2]~q ),
	.prn(vcc));
defparam \wr_addr[2] .is_wysiwyg = "true";
defparam \wr_addr[2] .power_up = "low";

dffeas \wr_addr[3] (
	.clk(clk),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\wr_addr[3]~q ),
	.prn(vcc));
defparam \wr_addr[3] .is_wysiwyg = "true";
defparam \wr_addr[3] .power_up = "low";

cyclonev_lcell_comb \Mux1~1 (
	.dataa(!\sw[0]~q ),
	.datab(!\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~1 .extended_lut = "off";
defparam \Mux1~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Mux1~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~2 (
	.dataa(!\sw[0]~q ),
	.datab(!\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~2 .extended_lut = "off";
defparam \Mux1~2 .lut_mask = 64'h7777777777777777;
defparam \Mux1~2 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!\sw[0]~q ),
	.datab(!\sw[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \anb~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!anb1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\anb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \anb~0 .extended_lut = "off";
defparam \anb~0 .lut_mask = 64'h6666666666666666;
defparam \anb~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_lpp_serial (
	data_real_o_0,
	data_real_o_1,
	data_real_o_2,
	data_real_o_3,
	data_real_o_4,
	data_real_o_5,
	data_real_o_6,
	data_real_o_7,
	tdl_arr_4,
	global_clock_enable,
	data_imag_o_0,
	data_imag_o_1,
	data_imag_o_2,
	data_imag_o_3,
	data_imag_o_4,
	data_imag_o_5,
	data_imag_o_6,
	data_imag_o_7,
	ram_in_reg_2_3,
	ram_in_reg_2_7,
	ram_in_reg_2_1,
	ram_in_reg_2_5,
	data_3_real_i,
	data_1_real_i,
	data_3_imag_i,
	data_1_imag_i,
	ram_in_reg_3_3,
	ram_in_reg_3_7,
	ram_in_reg_3_1,
	ram_in_reg_3_5,
	ram_in_reg_4_3,
	ram_in_reg_4_7,
	ram_in_reg_4_1,
	ram_in_reg_4_5,
	ram_in_reg_5_3,
	ram_in_reg_5_7,
	ram_in_reg_5_1,
	ram_in_reg_5_5,
	ram_in_reg_6_3,
	ram_in_reg_6_7,
	ram_in_reg_6_1,
	ram_in_reg_6_5,
	ram_in_reg_7_3,
	ram_in_reg_7_7,
	ram_in_reg_7_1,
	ram_in_reg_7_5,
	ram_in_reg_1_3,
	ram_in_reg_1_7,
	ram_in_reg_1_1,
	ram_in_reg_1_5,
	ram_in_reg_0_3,
	ram_in_reg_0_7,
	ram_in_reg_0_1,
	ram_in_reg_0_5,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	data_real_o_0;
output 	data_real_o_1;
output 	data_real_o_2;
output 	data_real_o_3;
output 	data_real_o_4;
output 	data_real_o_5;
output 	data_real_o_6;
output 	data_real_o_7;
input 	tdl_arr_4;
input 	global_clock_enable;
output 	data_imag_o_0;
output 	data_imag_o_1;
output 	data_imag_o_2;
output 	data_imag_o_3;
output 	data_imag_o_4;
output 	data_imag_o_5;
output 	data_imag_o_6;
output 	data_imag_o_7;
input 	ram_in_reg_2_3;
input 	ram_in_reg_2_7;
input 	ram_in_reg_2_1;
input 	ram_in_reg_2_5;
input 	[7:0] data_3_real_i;
input 	[7:0] data_1_real_i;
input 	[7:0] data_3_imag_i;
input 	[7:0] data_1_imag_i;
input 	ram_in_reg_3_3;
input 	ram_in_reg_3_7;
input 	ram_in_reg_3_1;
input 	ram_in_reg_3_5;
input 	ram_in_reg_4_3;
input 	ram_in_reg_4_7;
input 	ram_in_reg_4_1;
input 	ram_in_reg_4_5;
input 	ram_in_reg_5_3;
input 	ram_in_reg_5_7;
input 	ram_in_reg_5_1;
input 	ram_in_reg_5_5;
input 	ram_in_reg_6_3;
input 	ram_in_reg_6_7;
input 	ram_in_reg_6_1;
input 	ram_in_reg_6_5;
input 	ram_in_reg_7_3;
input 	ram_in_reg_7_7;
input 	ram_in_reg_7_1;
input 	ram_in_reg_7_5;
input 	ram_in_reg_1_3;
input 	ram_in_reg_1_7;
input 	ram_in_reg_1_1;
input 	ram_in_reg_1_5;
input 	ram_in_reg_0_3;
input 	ram_in_reg_0_7;
input 	ram_in_reg_0_1;
input 	ram_in_reg_0_5;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add9~1_sumout ;
wire \Add9~2 ;
wire \Add11~1_sumout ;
wire \Add11~2 ;
wire \Add9~5_sumout ;
wire \Add9~6 ;
wire \Add11~5_sumout ;
wire \Add11~6 ;
wire \Add9~9_sumout ;
wire \Add9~10 ;
wire \Add11~9_sumout ;
wire \Add11~10 ;
wire \Add9~13_sumout ;
wire \Add9~14 ;
wire \Add11~13_sumout ;
wire \Add11~14 ;
wire \Add9~17_sumout ;
wire \Add9~18 ;
wire \Add11~17_sumout ;
wire \Add11~18 ;
wire \Add9~21_sumout ;
wire \Add9~22 ;
wire \Add11~21_sumout ;
wire \Add11~22 ;
wire \Add9~25_sumout ;
wire \Add9~26 ;
wire \Add11~25_sumout ;
wire \Add11~26 ;
wire \Add9~29_sumout ;
wire \Add11~29_sumout ;
wire \Add9~33_sumout ;
wire \Add9~34 ;
wire \Add11~33_sumout ;
wire \Add11~34 ;
wire \Add3~1_sumout ;
wire \Add3~2 ;
wire \Add1~1_sumout ;
wire \Add1~2 ;
wire \Add9~37_sumout ;
wire \Add9~38 ;
wire \Add4~1_sumout ;
wire \Add4~2 ;
wire \Add2~1_sumout ;
wire \Add2~2 ;
wire \Add11~37_sumout ;
wire \Add11~38 ;
wire \Add3~5_sumout ;
wire \Add3~6 ;
wire \Add1~5_sumout ;
wire \Add1~6 ;
wire \Add4~5_sumout ;
wire \Add4~6 ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add3~9_sumout ;
wire \Add3~10 ;
wire \Add1~9_sumout ;
wire \Add1~10 ;
wire \Add4~9_sumout ;
wire \Add4~10 ;
wire \Add2~9_sumout ;
wire \Add2~10 ;
wire \Add3~13_sumout ;
wire \Add3~14 ;
wire \Add1~13_sumout ;
wire \Add1~14 ;
wire \Add4~13_sumout ;
wire \Add4~14 ;
wire \Add2~13_sumout ;
wire \Add2~14 ;
wire \Add3~17_sumout ;
wire \Add3~18 ;
wire \Add1~17_sumout ;
wire \Add1~18 ;
wire \Add4~17_sumout ;
wire \Add4~18 ;
wire \Add2~17_sumout ;
wire \Add2~18 ;
wire \Add3~21_sumout ;
wire \Add3~22 ;
wire \Add1~21_sumout ;
wire \Add1~22 ;
wire \Add4~21_sumout ;
wire \Add4~22 ;
wire \Add2~21_sumout ;
wire \Add2~22 ;
wire \Add3~25_sumout ;
wire \Add1~25_sumout ;
wire \Add4~25_sumout ;
wire \Add2~25_sumout ;
wire \add_in_r_d[2]~q ;
wire \add_in_r_c[2]~q ;
wire \Add3~29_sumout ;
wire \Add3~30 ;
wire \Add1~29_sumout ;
wire \Add1~30 ;
wire \Add9~42_cout ;
wire \add_in_i_d[2]~q ;
wire \add_in_i_c[2]~q ;
wire \Add4~29_sumout ;
wire \Add4~30 ;
wire \Add2~29_sumout ;
wire \Add2~30 ;
wire \Add11~42_cout ;
wire \add_in_r_d[3]~q ;
wire \add_in_r_c[3]~q ;
wire \add_in_i_d[3]~q ;
wire \add_in_i_c[3]~q ;
wire \add_in_r_d[4]~q ;
wire \add_in_r_c[4]~q ;
wire \add_in_i_d[4]~q ;
wire \add_in_i_c[4]~q ;
wire \add_in_r_d[5]~q ;
wire \add_in_r_c[5]~q ;
wire \add_in_i_d[5]~q ;
wire \add_in_i_c[5]~q ;
wire \add_in_r_d[6]~q ;
wire \add_in_r_c[6]~q ;
wire \add_in_i_d[6]~q ;
wire \add_in_i_c[6]~q ;
wire \add_in_r_d[7]~q ;
wire \add_in_r_c[7]~q ;
wire \add_in_i_d[7]~q ;
wire \add_in_i_c[7]~q ;
wire \add_in_r_d[1]~q ;
wire \add_in_r_c[1]~q ;
wire \Add3~33_sumout ;
wire \Add3~34 ;
wire \Add1~33_sumout ;
wire \Add1~34 ;
wire \add_in_i_d[1]~q ;
wire \add_in_i_c[1]~q ;
wire \Add4~33_sumout ;
wire \Add4~34 ;
wire \Add2~33_sumout ;
wire \Add2~34 ;
wire \add_in_r_d[0]~q ;
wire \add_in_r_c[0]~q ;
wire \Add3~38_cout ;
wire \Add1~38_cout ;
wire \add_in_i_d[0]~q ;
wire \add_in_i_c[0]~q ;
wire \Add4~38_cout ;
wire \Add2~38_cout ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \output_r[2]~q ;
wire \output_i[2]~q ;
wire \output_r[3]~q ;
wire \output_i[3]~q ;
wire \output_r[4]~q ;
wire \output_i[4]~q ;
wire \output_r[5]~q ;
wire \output_i[5]~q ;
wire \output_r[6]~q ;
wire \output_i[6]~q ;
wire \output_r[7]~q ;
wire \output_i[7]~q ;
wire \output_r[8]~q ;
wire \output_i[8]~q ;
wire \output_r[9]~q ;
wire \output_i[9]~q ;
wire \output_r[1]~q ;
wire \output_i[1]~q ;
wire \sgn_2r~q ;
wire \result_rb[2]~q ;
wire \result_ra[2]~q ;
wire \output_r[0]~q ;
wire \sgn_2i~q ;
wire \result_ib[2]~q ;
wire \result_ia[2]~q ;
wire \output_i[0]~q ;
wire \result_rb[3]~q ;
wire \result_ra[3]~q ;
wire \result_ib[3]~q ;
wire \result_ia[3]~q ;
wire \result_rb[4]~q ;
wire \result_ra[4]~q ;
wire \result_ib[4]~q ;
wire \result_ia[4]~q ;
wire \result_rb[5]~q ;
wire \result_ra[5]~q ;
wire \result_ib[5]~q ;
wire \result_ia[5]~q ;
wire \result_rb[6]~q ;
wire \result_ra[6]~q ;
wire \result_ib[6]~q ;
wire \result_ia[6]~q ;
wire \result_rb[7]~q ;
wire \result_ra[7]~q ;
wire \result_ib[7]~q ;
wire \result_ia[7]~q ;
wire \result_rb[8]~q ;
wire \result_ra[8]~q ;
wire \result_ib[8]~q ;
wire \result_ia[8]~q ;
wire \sign_vec[1]~q ;
wire \result_rb[1]~q ;
wire \result_ra[1]~q ;
wire \sign_vec[0]~q ;
wire \result_ib[1]~q ;
wire \result_ia[1]~q ;
wire \sign_sel[1]~q ;
wire \sign_vec[3]~q ;
wire \add_in_r_b[2]~q ;
wire \add_in_r_a[2]~q ;
wire \result_rb[0]~q ;
wire \result_ra[0]~q ;
wire \sign_sel[0]~q ;
wire \Mux0~0_combout ;
wire \add_in_i_b[2]~q ;
wire \add_in_i_a[2]~q ;
wire \result_ib[0]~q ;
wire \result_ia[0]~q ;
wire \add_in_r_b[3]~q ;
wire \add_in_r_a[3]~q ;
wire \add_in_i_b[3]~q ;
wire \add_in_i_a[3]~q ;
wire \add_in_r_b[4]~q ;
wire \add_in_r_a[4]~q ;
wire \add_in_i_b[4]~q ;
wire \add_in_i_a[4]~q ;
wire \add_in_r_b[5]~q ;
wire \add_in_r_a[5]~q ;
wire \add_in_i_b[5]~q ;
wire \add_in_i_a[5]~q ;
wire \add_in_r_b[6]~q ;
wire \add_in_r_a[6]~q ;
wire \add_in_i_b[6]~q ;
wire \add_in_i_a[6]~q ;
wire \add_in_r_b[7]~q ;
wire \add_in_r_a[7]~q ;
wire \add_in_i_b[7]~q ;
wire \add_in_i_a[7]~q ;
wire \offset_counter[5]~q ;
wire \add_in_r_b[1]~q ;
wire \add_in_r_a[1]~q ;
wire \offset_counter[4]~q ;
wire \add_in_i_b[1]~q ;
wire \add_in_i_a[1]~q ;
wire \offset_counter[3]~q ;
wire \offset_counter[2]~q ;
wire \offset_counter[0]~q ;
wire \offset_counter[1]~q ;
wire \Add0~0_combout ;
wire \offset_counter~0_combout ;
wire \add_in_r_b[0]~q ;
wire \add_in_r_a[0]~q ;
wire \offset_counter~1_combout ;
wire \add_in_i_b[0]~q ;
wire \add_in_i_a[0]~q ;
wire \offset_counter~2_combout ;
wire \offset_counter~3_combout ;
wire \offset_counter~4_combout ;
wire \offset_counter~5_combout ;
wire \sign_vec[1]~0_combout ;
wire \sign_vec[3]~2_combout ;
wire \data_imag_o[0]~0_combout ;
wire \data_imag_o[1]~1_combout ;
wire \data_imag_o[2]~2_combout ;
wire \data_imag_o[3]~3_combout ;
wire \data_imag_o[4]~4_combout ;
wire \data_imag_o[5]~5_combout ;
wire \data_imag_o[6]~6_combout ;
wire \data_imag_o[7]~7_combout ;


IFFT_asj_fft_pround_15 \gen_full_rnd:u1 (
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.output_i_2(\output_i[2]~q ),
	.output_i_3(\output_i[3]~q ),
	.output_i_4(\output_i[4]~q ),
	.output_i_5(\output_i[5]~q ),
	.output_i_6(\output_i[6]~q ),
	.output_i_7(\output_i[7]~q ),
	.output_i_8(\output_i[8]~q ),
	.output_i_9(\output_i[9]~q ),
	.output_i_1(\output_i[1]~q ),
	.output_i_0(\output_i[0]~q ),
	.clk(clk));

IFFT_asj_fft_pround_14 \gen_full_rnd:u0 (
	.global_clock_enable(global_clock_enable),
	.pipeline_dffe_2(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.output_r_2(\output_r[2]~q ),
	.output_r_3(\output_r[3]~q ),
	.output_r_4(\output_r[4]~q ),
	.output_r_5(\output_r[5]~q ),
	.output_r_6(\output_r[6]~q ),
	.output_r_7(\output_r[7]~q ),
	.output_r_8(\output_r[8]~q ),
	.output_r_9(\output_r[9]~q ),
	.output_r_1(\output_r[1]~q ),
	.output_r_0(\output_r[0]~q ),
	.clk(clk));

cyclonev_lcell_comb \Add9~1 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[2]~q ),
	.datae(gnd),
	.dataf(!\result_ra[2]~q ),
	.datag(gnd),
	.cin(\Add9~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~1_sumout ),
	.cout(\Add9~2 ),
	.shareout());
defparam \Add9~1 .extended_lut = "off";
defparam \Add9~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~1 .shared_arith = "off";

cyclonev_lcell_comb \Add11~1 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[2]~q ),
	.datae(gnd),
	.dataf(!\result_ia[2]~q ),
	.datag(gnd),
	.cin(\Add11~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~1_sumout ),
	.cout(\Add11~2 ),
	.shareout());
defparam \Add11~1 .extended_lut = "off";
defparam \Add11~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~1 .shared_arith = "off";

cyclonev_lcell_comb \Add9~5 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[3]~q ),
	.datae(gnd),
	.dataf(!\result_ra[3]~q ),
	.datag(gnd),
	.cin(\Add9~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~5_sumout ),
	.cout(\Add9~6 ),
	.shareout());
defparam \Add9~5 .extended_lut = "off";
defparam \Add9~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~5 .shared_arith = "off";

cyclonev_lcell_comb \Add11~5 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[3]~q ),
	.datae(gnd),
	.dataf(!\result_ia[3]~q ),
	.datag(gnd),
	.cin(\Add11~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~5_sumout ),
	.cout(\Add11~6 ),
	.shareout());
defparam \Add11~5 .extended_lut = "off";
defparam \Add11~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~5 .shared_arith = "off";

cyclonev_lcell_comb \Add9~9 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[4]~q ),
	.datae(gnd),
	.dataf(!\result_ra[4]~q ),
	.datag(gnd),
	.cin(\Add9~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~9_sumout ),
	.cout(\Add9~10 ),
	.shareout());
defparam \Add9~9 .extended_lut = "off";
defparam \Add9~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~9 .shared_arith = "off";

cyclonev_lcell_comb \Add11~9 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[4]~q ),
	.datae(gnd),
	.dataf(!\result_ia[4]~q ),
	.datag(gnd),
	.cin(\Add11~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~9_sumout ),
	.cout(\Add11~10 ),
	.shareout());
defparam \Add11~9 .extended_lut = "off";
defparam \Add11~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~9 .shared_arith = "off";

cyclonev_lcell_comb \Add9~13 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[5]~q ),
	.datae(gnd),
	.dataf(!\result_ra[5]~q ),
	.datag(gnd),
	.cin(\Add9~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~13_sumout ),
	.cout(\Add9~14 ),
	.shareout());
defparam \Add9~13 .extended_lut = "off";
defparam \Add9~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~13 .shared_arith = "off";

cyclonev_lcell_comb \Add11~13 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[5]~q ),
	.datae(gnd),
	.dataf(!\result_ia[5]~q ),
	.datag(gnd),
	.cin(\Add11~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~13_sumout ),
	.cout(\Add11~14 ),
	.shareout());
defparam \Add11~13 .extended_lut = "off";
defparam \Add11~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~13 .shared_arith = "off";

cyclonev_lcell_comb \Add9~17 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[6]~q ),
	.datae(gnd),
	.dataf(!\result_ra[6]~q ),
	.datag(gnd),
	.cin(\Add9~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~17_sumout ),
	.cout(\Add9~18 ),
	.shareout());
defparam \Add9~17 .extended_lut = "off";
defparam \Add9~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~17 .shared_arith = "off";

cyclonev_lcell_comb \Add11~17 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[6]~q ),
	.datae(gnd),
	.dataf(!\result_ia[6]~q ),
	.datag(gnd),
	.cin(\Add11~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~17_sumout ),
	.cout(\Add11~18 ),
	.shareout());
defparam \Add11~17 .extended_lut = "off";
defparam \Add11~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~17 .shared_arith = "off";

cyclonev_lcell_comb \Add9~21 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[7]~q ),
	.datae(gnd),
	.dataf(!\result_ra[7]~q ),
	.datag(gnd),
	.cin(\Add9~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~21_sumout ),
	.cout(\Add9~22 ),
	.shareout());
defparam \Add9~21 .extended_lut = "off";
defparam \Add9~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~21 .shared_arith = "off";

cyclonev_lcell_comb \Add11~21 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[7]~q ),
	.datae(gnd),
	.dataf(!\result_ia[7]~q ),
	.datag(gnd),
	.cin(\Add11~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~21_sumout ),
	.cout(\Add11~22 ),
	.shareout());
defparam \Add11~21 .extended_lut = "off";
defparam \Add11~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~21 .shared_arith = "off";

cyclonev_lcell_comb \Add9~25 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[8]~q ),
	.datae(gnd),
	.dataf(!\result_ra[8]~q ),
	.datag(gnd),
	.cin(\Add9~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~25_sumout ),
	.cout(\Add9~26 ),
	.shareout());
defparam \Add9~25 .extended_lut = "off";
defparam \Add9~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~25 .shared_arith = "off";

cyclonev_lcell_comb \Add11~25 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[8]~q ),
	.datae(gnd),
	.dataf(!\result_ia[8]~q ),
	.datag(gnd),
	.cin(\Add11~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~25_sumout ),
	.cout(\Add11~26 ),
	.shareout());
defparam \Add11~25 .extended_lut = "off";
defparam \Add11~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~25 .shared_arith = "off";

cyclonev_lcell_comb \Add9~29 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[8]~q ),
	.datae(gnd),
	.dataf(!\result_ra[8]~q ),
	.datag(gnd),
	.cin(\Add9~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~29_sumout ),
	.cout(),
	.shareout());
defparam \Add9~29 .extended_lut = "off";
defparam \Add9~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~29 .shared_arith = "off";

cyclonev_lcell_comb \Add11~29 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[8]~q ),
	.datae(gnd),
	.dataf(!\result_ia[8]~q ),
	.datag(gnd),
	.cin(\Add11~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~29_sumout ),
	.cout(),
	.shareout());
defparam \Add11~29 .extended_lut = "off";
defparam \Add11~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~29 .shared_arith = "off";

cyclonev_lcell_comb \Add9~33 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[1]~q ),
	.datae(gnd),
	.dataf(!\result_ra[1]~q ),
	.datag(gnd),
	.cin(\Add9~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~33_sumout ),
	.cout(\Add9~34 ),
	.shareout());
defparam \Add9~33 .extended_lut = "off";
defparam \Add9~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~33 .shared_arith = "off";

cyclonev_lcell_comb \Add11~33 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[1]~q ),
	.datae(gnd),
	.dataf(!\result_ia[1]~q ),
	.datag(gnd),
	.cin(\Add11~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~33_sumout ),
	.cout(\Add11~34 ),
	.shareout());
defparam \Add11~33 .extended_lut = "off";
defparam \Add11~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~33 .shared_arith = "off";

cyclonev_lcell_comb \Add3~1 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[2]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[2]~q ),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[2]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[2]~q ),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add9~37 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_rb[0]~q ),
	.datae(gnd),
	.dataf(!\result_ra[0]~q ),
	.datag(gnd),
	.cin(\Add9~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~37_sumout ),
	.cout(\Add9~38 ),
	.shareout());
defparam \Add9~37 .extended_lut = "off";
defparam \Add9~37 .lut_mask = 64'h0000FF00000055AA;
defparam \Add9~37 .shared_arith = "off";

cyclonev_lcell_comb \Add4~1 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[2]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[2]~q ),
	.datag(gnd),
	.cin(\Add4~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[2]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[2]~q ),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Add11~37 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\result_ib[0]~q ),
	.datae(gnd),
	.dataf(!\result_ia[0]~q ),
	.datag(gnd),
	.cin(\Add11~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~37_sumout ),
	.cout(\Add11~38 ),
	.shareout());
defparam \Add11~37 .extended_lut = "off";
defparam \Add11~37 .lut_mask = 64'h0000FF00000055AA;
defparam \Add11~37 .shared_arith = "off";

cyclonev_lcell_comb \Add3~5 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[3]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[3]~q ),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[3]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[3]~q ),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[3]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[3]~q ),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add2~5 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[3]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[3]~q ),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \Add3~9 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[4]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[4]~q ),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[4]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[4]~q ),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[4]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[4]~q ),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add2~9 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[4]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[4]~q ),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \Add3~13 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[5]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[5]~q ),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[5]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[5]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[5]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[5]~q ),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add2~13 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[5]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[5]~q ),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \Add3~17 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[6]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[6]~q ),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[6]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[6]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[6]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[6]~q ),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add2~17 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[6]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[6]~q ),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~17 .shared_arith = "off";

cyclonev_lcell_comb \Add3~21 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[7]~q ),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[7]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add4~21 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[7]~q ),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(\Add4~22 ),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~21 .shared_arith = "off";

cyclonev_lcell_comb \Add2~21 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[7]~q ),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~21 .shared_arith = "off";

cyclonev_lcell_comb \Add3~25 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[7]~q ),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[7]~q ),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[7]~q ),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(),
	.shareout());
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~25 .shared_arith = "off";

cyclonev_lcell_comb \Add2~25 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[7]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[7]~q ),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(),
	.shareout());
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~25 .shared_arith = "off";

dffeas \add_in_r_d[2] (
	.clk(clk),
	.d(ram_in_reg_2_3),
	.asdata(ram_in_reg_2_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[2]~q ),
	.prn(vcc));
defparam \add_in_r_d[2] .is_wysiwyg = "true";
defparam \add_in_r_d[2] .power_up = "low";

dffeas \add_in_r_c[2] (
	.clk(clk),
	.d(ram_in_reg_2_1),
	.asdata(ram_in_reg_2_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[2]~q ),
	.prn(vcc));
defparam \add_in_r_c[2] .is_wysiwyg = "true";
defparam \add_in_r_c[2] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[1]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[1]~q ),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[1]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[1]~q ),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~29 .shared_arith = "off";

cyclonev_lcell_comb \Add9~42 (
	.dataa(!\sgn_2r~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add9~42_cout ),
	.shareout());
defparam \Add9~42 .extended_lut = "off";
defparam \Add9~42 .lut_mask = 64'h000000000000AAAA;
defparam \Add9~42 .shared_arith = "off";

dffeas \add_in_i_d[2] (
	.clk(clk),
	.d(ram_in_reg_2_7),
	.asdata(ram_in_reg_2_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[2]~q ),
	.prn(vcc));
defparam \add_in_i_d[2] .is_wysiwyg = "true";
defparam \add_in_i_d[2] .power_up = "low";

dffeas \add_in_i_c[2] (
	.clk(clk),
	.d(ram_in_reg_2_5),
	.asdata(ram_in_reg_2_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[2]~q ),
	.prn(vcc));
defparam \add_in_i_c[2] .is_wysiwyg = "true";
defparam \add_in_i_c[2] .power_up = "low";

cyclonev_lcell_comb \Add4~29 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[1]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[1]~q ),
	.datag(gnd),
	.cin(\Add4~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~29_sumout ),
	.cout(\Add4~30 ),
	.shareout());
defparam \Add4~29 .extended_lut = "off";
defparam \Add4~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~29 .shared_arith = "off";

cyclonev_lcell_comb \Add2~29 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[1]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[1]~q ),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout());
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~29 .shared_arith = "off";

cyclonev_lcell_comb \Add11~42 (
	.dataa(!\sgn_2i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add11~42_cout ),
	.shareout());
defparam \Add11~42 .extended_lut = "off";
defparam \Add11~42 .lut_mask = 64'h000000000000AAAA;
defparam \Add11~42 .shared_arith = "off";

dffeas \add_in_r_d[3] (
	.clk(clk),
	.d(ram_in_reg_3_3),
	.asdata(ram_in_reg_3_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[3]~q ),
	.prn(vcc));
defparam \add_in_r_d[3] .is_wysiwyg = "true";
defparam \add_in_r_d[3] .power_up = "low";

dffeas \add_in_r_c[3] (
	.clk(clk),
	.d(ram_in_reg_3_1),
	.asdata(ram_in_reg_3_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[3]~q ),
	.prn(vcc));
defparam \add_in_r_c[3] .is_wysiwyg = "true";
defparam \add_in_r_c[3] .power_up = "low";

dffeas \add_in_i_d[3] (
	.clk(clk),
	.d(ram_in_reg_3_7),
	.asdata(ram_in_reg_3_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[3]~q ),
	.prn(vcc));
defparam \add_in_i_d[3] .is_wysiwyg = "true";
defparam \add_in_i_d[3] .power_up = "low";

dffeas \add_in_i_c[3] (
	.clk(clk),
	.d(ram_in_reg_3_5),
	.asdata(ram_in_reg_3_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[3]~q ),
	.prn(vcc));
defparam \add_in_i_c[3] .is_wysiwyg = "true";
defparam \add_in_i_c[3] .power_up = "low";

dffeas \add_in_r_d[4] (
	.clk(clk),
	.d(ram_in_reg_4_3),
	.asdata(ram_in_reg_4_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[4]~q ),
	.prn(vcc));
defparam \add_in_r_d[4] .is_wysiwyg = "true";
defparam \add_in_r_d[4] .power_up = "low";

dffeas \add_in_r_c[4] (
	.clk(clk),
	.d(ram_in_reg_4_1),
	.asdata(ram_in_reg_4_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[4]~q ),
	.prn(vcc));
defparam \add_in_r_c[4] .is_wysiwyg = "true";
defparam \add_in_r_c[4] .power_up = "low";

dffeas \add_in_i_d[4] (
	.clk(clk),
	.d(ram_in_reg_4_7),
	.asdata(ram_in_reg_4_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[4]~q ),
	.prn(vcc));
defparam \add_in_i_d[4] .is_wysiwyg = "true";
defparam \add_in_i_d[4] .power_up = "low";

dffeas \add_in_i_c[4] (
	.clk(clk),
	.d(ram_in_reg_4_5),
	.asdata(ram_in_reg_4_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[4]~q ),
	.prn(vcc));
defparam \add_in_i_c[4] .is_wysiwyg = "true";
defparam \add_in_i_c[4] .power_up = "low";

dffeas \add_in_r_d[5] (
	.clk(clk),
	.d(ram_in_reg_5_3),
	.asdata(ram_in_reg_5_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[5]~q ),
	.prn(vcc));
defparam \add_in_r_d[5] .is_wysiwyg = "true";
defparam \add_in_r_d[5] .power_up = "low";

dffeas \add_in_r_c[5] (
	.clk(clk),
	.d(ram_in_reg_5_1),
	.asdata(ram_in_reg_5_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[5]~q ),
	.prn(vcc));
defparam \add_in_r_c[5] .is_wysiwyg = "true";
defparam \add_in_r_c[5] .power_up = "low";

dffeas \add_in_i_d[5] (
	.clk(clk),
	.d(ram_in_reg_5_7),
	.asdata(ram_in_reg_5_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[5]~q ),
	.prn(vcc));
defparam \add_in_i_d[5] .is_wysiwyg = "true";
defparam \add_in_i_d[5] .power_up = "low";

dffeas \add_in_i_c[5] (
	.clk(clk),
	.d(ram_in_reg_5_5),
	.asdata(ram_in_reg_5_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[5]~q ),
	.prn(vcc));
defparam \add_in_i_c[5] .is_wysiwyg = "true";
defparam \add_in_i_c[5] .power_up = "low";

dffeas \add_in_r_d[6] (
	.clk(clk),
	.d(ram_in_reg_6_3),
	.asdata(ram_in_reg_6_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[6]~q ),
	.prn(vcc));
defparam \add_in_r_d[6] .is_wysiwyg = "true";
defparam \add_in_r_d[6] .power_up = "low";

dffeas \add_in_r_c[6] (
	.clk(clk),
	.d(ram_in_reg_6_1),
	.asdata(ram_in_reg_6_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[6]~q ),
	.prn(vcc));
defparam \add_in_r_c[6] .is_wysiwyg = "true";
defparam \add_in_r_c[6] .power_up = "low";

dffeas \add_in_i_d[6] (
	.clk(clk),
	.d(ram_in_reg_6_7),
	.asdata(ram_in_reg_6_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[6]~q ),
	.prn(vcc));
defparam \add_in_i_d[6] .is_wysiwyg = "true";
defparam \add_in_i_d[6] .power_up = "low";

dffeas \add_in_i_c[6] (
	.clk(clk),
	.d(ram_in_reg_6_5),
	.asdata(ram_in_reg_6_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[6]~q ),
	.prn(vcc));
defparam \add_in_i_c[6] .is_wysiwyg = "true";
defparam \add_in_i_c[6] .power_up = "low";

dffeas \add_in_r_d[7] (
	.clk(clk),
	.d(ram_in_reg_7_3),
	.asdata(ram_in_reg_7_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[7]~q ),
	.prn(vcc));
defparam \add_in_r_d[7] .is_wysiwyg = "true";
defparam \add_in_r_d[7] .power_up = "low";

dffeas \add_in_r_c[7] (
	.clk(clk),
	.d(ram_in_reg_7_1),
	.asdata(ram_in_reg_7_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[7]~q ),
	.prn(vcc));
defparam \add_in_r_c[7] .is_wysiwyg = "true";
defparam \add_in_r_c[7] .power_up = "low";

dffeas \add_in_i_d[7] (
	.clk(clk),
	.d(ram_in_reg_7_7),
	.asdata(ram_in_reg_7_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[7]~q ),
	.prn(vcc));
defparam \add_in_i_d[7] .is_wysiwyg = "true";
defparam \add_in_i_d[7] .power_up = "low";

dffeas \add_in_i_c[7] (
	.clk(clk),
	.d(ram_in_reg_7_5),
	.asdata(ram_in_reg_7_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[7]~q ),
	.prn(vcc));
defparam \add_in_i_c[7] .is_wysiwyg = "true";
defparam \add_in_i_c[7] .power_up = "low";

dffeas \add_in_r_d[1] (
	.clk(clk),
	.d(ram_in_reg_1_3),
	.asdata(ram_in_reg_1_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[1]~q ),
	.prn(vcc));
defparam \add_in_r_d[1] .is_wysiwyg = "true";
defparam \add_in_r_d[1] .power_up = "low";

dffeas \add_in_r_c[1] (
	.clk(clk),
	.d(ram_in_reg_1_1),
	.asdata(ram_in_reg_1_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[1]~q ),
	.prn(vcc));
defparam \add_in_r_c[1] .is_wysiwyg = "true";
defparam \add_in_r_c[1] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_d[0]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_c[0]~q ),
	.datag(gnd),
	.cin(\Add3~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add3~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_r_b[0]~q ),
	.datae(gnd),
	.dataf(!\add_in_r_a[0]~q ),
	.datag(gnd),
	.cin(\Add1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add1~33 .shared_arith = "off";

dffeas \add_in_i_d[1] (
	.clk(clk),
	.d(ram_in_reg_1_7),
	.asdata(ram_in_reg_1_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[1]~q ),
	.prn(vcc));
defparam \add_in_i_d[1] .is_wysiwyg = "true";
defparam \add_in_i_d[1] .power_up = "low";

dffeas \add_in_i_c[1] (
	.clk(clk),
	.d(ram_in_reg_1_5),
	.asdata(ram_in_reg_1_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[1]~q ),
	.prn(vcc));
defparam \add_in_i_c[1] .is_wysiwyg = "true";
defparam \add_in_i_c[1] .power_up = "low";

cyclonev_lcell_comb \Add4~33 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_d[0]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_c[0]~q ),
	.datag(gnd),
	.cin(\Add4~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~33_sumout ),
	.cout(\Add4~34 ),
	.shareout());
defparam \Add4~33 .extended_lut = "off";
defparam \Add4~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add4~33 .shared_arith = "off";

cyclonev_lcell_comb \Add2~33 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\add_in_i_b[0]~q ),
	.datae(gnd),
	.dataf(!\add_in_i_a[0]~q ),
	.datag(gnd),
	.cin(\Add2~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout());
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add2~33 .shared_arith = "off";

dffeas \add_in_r_d[0] (
	.clk(clk),
	.d(ram_in_reg_0_3),
	.asdata(ram_in_reg_0_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_d[0]~q ),
	.prn(vcc));
defparam \add_in_r_d[0] .is_wysiwyg = "true";
defparam \add_in_r_d[0] .power_up = "low";

dffeas \add_in_r_c[0] (
	.clk(clk),
	.d(ram_in_reg_0_1),
	.asdata(ram_in_reg_0_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_r_c[0]~q ),
	.prn(vcc));
defparam \add_in_r_c[0] .is_wysiwyg = "true";
defparam \add_in_r_c[0] .power_up = "low";

cyclonev_lcell_comb \Add3~38 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add3~38_cout ),
	.shareout());
defparam \Add3~38 .extended_lut = "off";
defparam \Add3~38 .lut_mask = 64'h000000000000AAAA;
defparam \Add3~38 .shared_arith = "off";

cyclonev_lcell_comb \Add1~38 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add1~38_cout ),
	.shareout());
defparam \Add1~38 .extended_lut = "off";
defparam \Add1~38 .lut_mask = 64'h000000000000AAAA;
defparam \Add1~38 .shared_arith = "off";

dffeas \add_in_i_d[0] (
	.clk(clk),
	.d(ram_in_reg_0_7),
	.asdata(ram_in_reg_0_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_d[0]~q ),
	.prn(vcc));
defparam \add_in_i_d[0] .is_wysiwyg = "true";
defparam \add_in_i_d[0] .power_up = "low";

dffeas \add_in_i_c[0] (
	.clk(clk),
	.d(ram_in_reg_0_5),
	.asdata(ram_in_reg_0_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sign_sel[0]~q ),
	.ena(!global_clock_enable),
	.q(\add_in_i_c[0]~q ),
	.prn(vcc));
defparam \add_in_i_c[0] .is_wysiwyg = "true";
defparam \add_in_i_c[0] .power_up = "low";

cyclonev_lcell_comb \Add4~38 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add4~38_cout ),
	.shareout());
defparam \Add4~38 .extended_lut = "off";
defparam \Add4~38 .lut_mask = 64'h000000000000AAAA;
defparam \Add4~38 .shared_arith = "off";

cyclonev_lcell_comb \Add2~38 (
	.dataa(!\sign_vec[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add2~38_cout ),
	.shareout());
defparam \Add2~38 .extended_lut = "off";
defparam \Add2~38 .lut_mask = 64'h000000000000AAAA;
defparam \Add2~38 .shared_arith = "off";

dffeas \output_r[2] (
	.clk(clk),
	.d(\Add9~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[2]~q ),
	.prn(vcc));
defparam \output_r[2] .is_wysiwyg = "true";
defparam \output_r[2] .power_up = "low";

dffeas \output_i[2] (
	.clk(clk),
	.d(\Add11~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[2]~q ),
	.prn(vcc));
defparam \output_i[2] .is_wysiwyg = "true";
defparam \output_i[2] .power_up = "low";

dffeas \output_r[3] (
	.clk(clk),
	.d(\Add9~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[3]~q ),
	.prn(vcc));
defparam \output_r[3] .is_wysiwyg = "true";
defparam \output_r[3] .power_up = "low";

dffeas \output_i[3] (
	.clk(clk),
	.d(\Add11~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[3]~q ),
	.prn(vcc));
defparam \output_i[3] .is_wysiwyg = "true";
defparam \output_i[3] .power_up = "low";

dffeas \output_r[4] (
	.clk(clk),
	.d(\Add9~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[4]~q ),
	.prn(vcc));
defparam \output_r[4] .is_wysiwyg = "true";
defparam \output_r[4] .power_up = "low";

dffeas \output_i[4] (
	.clk(clk),
	.d(\Add11~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[4]~q ),
	.prn(vcc));
defparam \output_i[4] .is_wysiwyg = "true";
defparam \output_i[4] .power_up = "low";

dffeas \output_r[5] (
	.clk(clk),
	.d(\Add9~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[5]~q ),
	.prn(vcc));
defparam \output_r[5] .is_wysiwyg = "true";
defparam \output_r[5] .power_up = "low";

dffeas \output_i[5] (
	.clk(clk),
	.d(\Add11~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[5]~q ),
	.prn(vcc));
defparam \output_i[5] .is_wysiwyg = "true";
defparam \output_i[5] .power_up = "low";

dffeas \output_r[6] (
	.clk(clk),
	.d(\Add9~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[6]~q ),
	.prn(vcc));
defparam \output_r[6] .is_wysiwyg = "true";
defparam \output_r[6] .power_up = "low";

dffeas \output_i[6] (
	.clk(clk),
	.d(\Add11~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[6]~q ),
	.prn(vcc));
defparam \output_i[6] .is_wysiwyg = "true";
defparam \output_i[6] .power_up = "low";

dffeas \output_r[7] (
	.clk(clk),
	.d(\Add9~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[7]~q ),
	.prn(vcc));
defparam \output_r[7] .is_wysiwyg = "true";
defparam \output_r[7] .power_up = "low";

dffeas \output_i[7] (
	.clk(clk),
	.d(\Add11~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[7]~q ),
	.prn(vcc));
defparam \output_i[7] .is_wysiwyg = "true";
defparam \output_i[7] .power_up = "low";

dffeas \output_r[8] (
	.clk(clk),
	.d(\Add9~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[8]~q ),
	.prn(vcc));
defparam \output_r[8] .is_wysiwyg = "true";
defparam \output_r[8] .power_up = "low";

dffeas \output_i[8] (
	.clk(clk),
	.d(\Add11~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[8]~q ),
	.prn(vcc));
defparam \output_i[8] .is_wysiwyg = "true";
defparam \output_i[8] .power_up = "low";

dffeas \output_r[9] (
	.clk(clk),
	.d(\Add9~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[9]~q ),
	.prn(vcc));
defparam \output_r[9] .is_wysiwyg = "true";
defparam \output_r[9] .power_up = "low";

dffeas \output_i[9] (
	.clk(clk),
	.d(\Add11~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[9]~q ),
	.prn(vcc));
defparam \output_i[9] .is_wysiwyg = "true";
defparam \output_i[9] .power_up = "low";

dffeas \output_r[1] (
	.clk(clk),
	.d(\Add9~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[1]~q ),
	.prn(vcc));
defparam \output_r[1] .is_wysiwyg = "true";
defparam \output_r[1] .power_up = "low";

dffeas \output_i[1] (
	.clk(clk),
	.d(\Add11~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[1]~q ),
	.prn(vcc));
defparam \output_i[1] .is_wysiwyg = "true";
defparam \output_i[1] .power_up = "low";

dffeas sgn_2r(
	.clk(clk),
	.d(\sign_vec[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sgn_2r~q ),
	.prn(vcc));
defparam sgn_2r.is_wysiwyg = "true";
defparam sgn_2r.power_up = "low";

dffeas \result_rb[2] (
	.clk(clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[2]~q ),
	.prn(vcc));
defparam \result_rb[2] .is_wysiwyg = "true";
defparam \result_rb[2] .power_up = "low";

dffeas \result_ra[2] (
	.clk(clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[2]~q ),
	.prn(vcc));
defparam \result_ra[2] .is_wysiwyg = "true";
defparam \result_ra[2] .power_up = "low";

dffeas \output_r[0] (
	.clk(clk),
	.d(\Add9~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_r[0]~q ),
	.prn(vcc));
defparam \output_r[0] .is_wysiwyg = "true";
defparam \output_r[0] .power_up = "low";

dffeas sgn_2i(
	.clk(clk),
	.d(\sign_vec[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sgn_2i~q ),
	.prn(vcc));
defparam sgn_2i.is_wysiwyg = "true";
defparam sgn_2i.power_up = "low";

dffeas \result_ib[2] (
	.clk(clk),
	.d(\Add4~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[2]~q ),
	.prn(vcc));
defparam \result_ib[2] .is_wysiwyg = "true";
defparam \result_ib[2] .power_up = "low";

dffeas \result_ia[2] (
	.clk(clk),
	.d(\Add2~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[2]~q ),
	.prn(vcc));
defparam \result_ia[2] .is_wysiwyg = "true";
defparam \result_ia[2] .power_up = "low";

dffeas \output_i[0] (
	.clk(clk),
	.d(\Add11~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\output_i[0]~q ),
	.prn(vcc));
defparam \output_i[0] .is_wysiwyg = "true";
defparam \output_i[0] .power_up = "low";

dffeas \result_rb[3] (
	.clk(clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[3]~q ),
	.prn(vcc));
defparam \result_rb[3] .is_wysiwyg = "true";
defparam \result_rb[3] .power_up = "low";

dffeas \result_ra[3] (
	.clk(clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[3]~q ),
	.prn(vcc));
defparam \result_ra[3] .is_wysiwyg = "true";
defparam \result_ra[3] .power_up = "low";

dffeas \result_ib[3] (
	.clk(clk),
	.d(\Add4~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[3]~q ),
	.prn(vcc));
defparam \result_ib[3] .is_wysiwyg = "true";
defparam \result_ib[3] .power_up = "low";

dffeas \result_ia[3] (
	.clk(clk),
	.d(\Add2~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[3]~q ),
	.prn(vcc));
defparam \result_ia[3] .is_wysiwyg = "true";
defparam \result_ia[3] .power_up = "low";

dffeas \result_rb[4] (
	.clk(clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[4]~q ),
	.prn(vcc));
defparam \result_rb[4] .is_wysiwyg = "true";
defparam \result_rb[4] .power_up = "low";

dffeas \result_ra[4] (
	.clk(clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[4]~q ),
	.prn(vcc));
defparam \result_ra[4] .is_wysiwyg = "true";
defparam \result_ra[4] .power_up = "low";

dffeas \result_ib[4] (
	.clk(clk),
	.d(\Add4~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[4]~q ),
	.prn(vcc));
defparam \result_ib[4] .is_wysiwyg = "true";
defparam \result_ib[4] .power_up = "low";

dffeas \result_ia[4] (
	.clk(clk),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[4]~q ),
	.prn(vcc));
defparam \result_ia[4] .is_wysiwyg = "true";
defparam \result_ia[4] .power_up = "low";

dffeas \result_rb[5] (
	.clk(clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[5]~q ),
	.prn(vcc));
defparam \result_rb[5] .is_wysiwyg = "true";
defparam \result_rb[5] .power_up = "low";

dffeas \result_ra[5] (
	.clk(clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[5]~q ),
	.prn(vcc));
defparam \result_ra[5] .is_wysiwyg = "true";
defparam \result_ra[5] .power_up = "low";

dffeas \result_ib[5] (
	.clk(clk),
	.d(\Add4~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[5]~q ),
	.prn(vcc));
defparam \result_ib[5] .is_wysiwyg = "true";
defparam \result_ib[5] .power_up = "low";

dffeas \result_ia[5] (
	.clk(clk),
	.d(\Add2~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[5]~q ),
	.prn(vcc));
defparam \result_ia[5] .is_wysiwyg = "true";
defparam \result_ia[5] .power_up = "low";

dffeas \result_rb[6] (
	.clk(clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[6]~q ),
	.prn(vcc));
defparam \result_rb[6] .is_wysiwyg = "true";
defparam \result_rb[6] .power_up = "low";

dffeas \result_ra[6] (
	.clk(clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[6]~q ),
	.prn(vcc));
defparam \result_ra[6] .is_wysiwyg = "true";
defparam \result_ra[6] .power_up = "low";

dffeas \result_ib[6] (
	.clk(clk),
	.d(\Add4~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[6]~q ),
	.prn(vcc));
defparam \result_ib[6] .is_wysiwyg = "true";
defparam \result_ib[6] .power_up = "low";

dffeas \result_ia[6] (
	.clk(clk),
	.d(\Add2~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[6]~q ),
	.prn(vcc));
defparam \result_ia[6] .is_wysiwyg = "true";
defparam \result_ia[6] .power_up = "low";

dffeas \result_rb[7] (
	.clk(clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[7]~q ),
	.prn(vcc));
defparam \result_rb[7] .is_wysiwyg = "true";
defparam \result_rb[7] .power_up = "low";

dffeas \result_ra[7] (
	.clk(clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[7]~q ),
	.prn(vcc));
defparam \result_ra[7] .is_wysiwyg = "true";
defparam \result_ra[7] .power_up = "low";

dffeas \result_ib[7] (
	.clk(clk),
	.d(\Add4~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[7]~q ),
	.prn(vcc));
defparam \result_ib[7] .is_wysiwyg = "true";
defparam \result_ib[7] .power_up = "low";

dffeas \result_ia[7] (
	.clk(clk),
	.d(\Add2~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[7]~q ),
	.prn(vcc));
defparam \result_ia[7] .is_wysiwyg = "true";
defparam \result_ia[7] .power_up = "low";

dffeas \result_rb[8] (
	.clk(clk),
	.d(\Add3~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[8]~q ),
	.prn(vcc));
defparam \result_rb[8] .is_wysiwyg = "true";
defparam \result_rb[8] .power_up = "low";

dffeas \result_ra[8] (
	.clk(clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[8]~q ),
	.prn(vcc));
defparam \result_ra[8] .is_wysiwyg = "true";
defparam \result_ra[8] .power_up = "low";

dffeas \result_ib[8] (
	.clk(clk),
	.d(\Add4~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[8]~q ),
	.prn(vcc));
defparam \result_ib[8] .is_wysiwyg = "true";
defparam \result_ib[8] .power_up = "low";

dffeas \result_ia[8] (
	.clk(clk),
	.d(\Add2~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[8]~q ),
	.prn(vcc));
defparam \result_ia[8] .is_wysiwyg = "true";
defparam \result_ia[8] .power_up = "low";

dffeas \sign_vec[1] (
	.clk(clk),
	.d(\sign_vec[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sign_vec[1]~q ),
	.prn(vcc));
defparam \sign_vec[1] .is_wysiwyg = "true";
defparam \sign_vec[1] .power_up = "low";

dffeas \result_rb[1] (
	.clk(clk),
	.d(\Add3~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[1]~q ),
	.prn(vcc));
defparam \result_rb[1] .is_wysiwyg = "true";
defparam \result_rb[1] .power_up = "low";

dffeas \result_ra[1] (
	.clk(clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[1]~q ),
	.prn(vcc));
defparam \result_ra[1] .is_wysiwyg = "true";
defparam \result_ra[1] .power_up = "low";

dffeas \sign_vec[0] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sign_vec[0]~q ),
	.prn(vcc));
defparam \sign_vec[0] .is_wysiwyg = "true";
defparam \sign_vec[0] .power_up = "low";

dffeas \result_ib[1] (
	.clk(clk),
	.d(\Add4~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[1]~q ),
	.prn(vcc));
defparam \result_ib[1] .is_wysiwyg = "true";
defparam \result_ib[1] .power_up = "low";

dffeas \result_ia[1] (
	.clk(clk),
	.d(\Add2~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[1]~q ),
	.prn(vcc));
defparam \result_ia[1] .is_wysiwyg = "true";
defparam \result_ia[1] .power_up = "low";

dffeas \sign_sel[1] (
	.clk(clk),
	.d(\offset_counter[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sign_sel[1]~q ),
	.prn(vcc));
defparam \sign_sel[1] .is_wysiwyg = "true";
defparam \sign_sel[1] .power_up = "low";

dffeas \sign_vec[3] (
	.clk(clk),
	.d(\sign_vec[3]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sign_vec[3]~q ),
	.prn(vcc));
defparam \sign_vec[3] .is_wysiwyg = "true";
defparam \sign_vec[3] .power_up = "low";

dffeas \add_in_r_b[2] (
	.clk(clk),
	.d(data_3_real_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[2]~q ),
	.prn(vcc));
defparam \add_in_r_b[2] .is_wysiwyg = "true";
defparam \add_in_r_b[2] .power_up = "low";

dffeas \add_in_r_a[2] (
	.clk(clk),
	.d(data_1_real_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[2]~q ),
	.prn(vcc));
defparam \add_in_r_a[2] .is_wysiwyg = "true";
defparam \add_in_r_a[2] .power_up = "low";

dffeas \result_rb[0] (
	.clk(clk),
	.d(\Add3~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_rb[0]~q ),
	.prn(vcc));
defparam \result_rb[0] .is_wysiwyg = "true";
defparam \result_rb[0] .power_up = "low";

dffeas \result_ra[0] (
	.clk(clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ra[0]~q ),
	.prn(vcc));
defparam \result_ra[0] .is_wysiwyg = "true";
defparam \result_ra[0] .power_up = "low";

dffeas \sign_sel[0] (
	.clk(clk),
	.d(\offset_counter[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\sign_sel[0]~q ),
	.prn(vcc));
defparam \sign_sel[0] .is_wysiwyg = "true";
defparam \sign_sel[0] .power_up = "low";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!\sign_sel[1]~q ),
	.datab(!\sign_sel[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h6666666666666666;
defparam \Mux0~0 .shared_arith = "off";

dffeas \add_in_i_b[2] (
	.clk(clk),
	.d(data_3_imag_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[2]~q ),
	.prn(vcc));
defparam \add_in_i_b[2] .is_wysiwyg = "true";
defparam \add_in_i_b[2] .power_up = "low";

dffeas \add_in_i_a[2] (
	.clk(clk),
	.d(data_1_imag_i[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[2]~q ),
	.prn(vcc));
defparam \add_in_i_a[2] .is_wysiwyg = "true";
defparam \add_in_i_a[2] .power_up = "low";

dffeas \result_ib[0] (
	.clk(clk),
	.d(\Add4~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ib[0]~q ),
	.prn(vcc));
defparam \result_ib[0] .is_wysiwyg = "true";
defparam \result_ib[0] .power_up = "low";

dffeas \result_ia[0] (
	.clk(clk),
	.d(\Add2~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\result_ia[0]~q ),
	.prn(vcc));
defparam \result_ia[0] .is_wysiwyg = "true";
defparam \result_ia[0] .power_up = "low";

dffeas \add_in_r_b[3] (
	.clk(clk),
	.d(data_3_real_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[3]~q ),
	.prn(vcc));
defparam \add_in_r_b[3] .is_wysiwyg = "true";
defparam \add_in_r_b[3] .power_up = "low";

dffeas \add_in_r_a[3] (
	.clk(clk),
	.d(data_1_real_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[3]~q ),
	.prn(vcc));
defparam \add_in_r_a[3] .is_wysiwyg = "true";
defparam \add_in_r_a[3] .power_up = "low";

dffeas \add_in_i_b[3] (
	.clk(clk),
	.d(data_3_imag_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[3]~q ),
	.prn(vcc));
defparam \add_in_i_b[3] .is_wysiwyg = "true";
defparam \add_in_i_b[3] .power_up = "low";

dffeas \add_in_i_a[3] (
	.clk(clk),
	.d(data_1_imag_i[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[3]~q ),
	.prn(vcc));
defparam \add_in_i_a[3] .is_wysiwyg = "true";
defparam \add_in_i_a[3] .power_up = "low";

dffeas \add_in_r_b[4] (
	.clk(clk),
	.d(data_3_real_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[4]~q ),
	.prn(vcc));
defparam \add_in_r_b[4] .is_wysiwyg = "true";
defparam \add_in_r_b[4] .power_up = "low";

dffeas \add_in_r_a[4] (
	.clk(clk),
	.d(data_1_real_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[4]~q ),
	.prn(vcc));
defparam \add_in_r_a[4] .is_wysiwyg = "true";
defparam \add_in_r_a[4] .power_up = "low";

dffeas \add_in_i_b[4] (
	.clk(clk),
	.d(data_3_imag_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[4]~q ),
	.prn(vcc));
defparam \add_in_i_b[4] .is_wysiwyg = "true";
defparam \add_in_i_b[4] .power_up = "low";

dffeas \add_in_i_a[4] (
	.clk(clk),
	.d(data_1_imag_i[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[4]~q ),
	.prn(vcc));
defparam \add_in_i_a[4] .is_wysiwyg = "true";
defparam \add_in_i_a[4] .power_up = "low";

dffeas \add_in_r_b[5] (
	.clk(clk),
	.d(data_3_real_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[5]~q ),
	.prn(vcc));
defparam \add_in_r_b[5] .is_wysiwyg = "true";
defparam \add_in_r_b[5] .power_up = "low";

dffeas \add_in_r_a[5] (
	.clk(clk),
	.d(data_1_real_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[5]~q ),
	.prn(vcc));
defparam \add_in_r_a[5] .is_wysiwyg = "true";
defparam \add_in_r_a[5] .power_up = "low";

dffeas \add_in_i_b[5] (
	.clk(clk),
	.d(data_3_imag_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[5]~q ),
	.prn(vcc));
defparam \add_in_i_b[5] .is_wysiwyg = "true";
defparam \add_in_i_b[5] .power_up = "low";

dffeas \add_in_i_a[5] (
	.clk(clk),
	.d(data_1_imag_i[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[5]~q ),
	.prn(vcc));
defparam \add_in_i_a[5] .is_wysiwyg = "true";
defparam \add_in_i_a[5] .power_up = "low";

dffeas \add_in_r_b[6] (
	.clk(clk),
	.d(data_3_real_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[6]~q ),
	.prn(vcc));
defparam \add_in_r_b[6] .is_wysiwyg = "true";
defparam \add_in_r_b[6] .power_up = "low";

dffeas \add_in_r_a[6] (
	.clk(clk),
	.d(data_1_real_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[6]~q ),
	.prn(vcc));
defparam \add_in_r_a[6] .is_wysiwyg = "true";
defparam \add_in_r_a[6] .power_up = "low";

dffeas \add_in_i_b[6] (
	.clk(clk),
	.d(data_3_imag_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[6]~q ),
	.prn(vcc));
defparam \add_in_i_b[6] .is_wysiwyg = "true";
defparam \add_in_i_b[6] .power_up = "low";

dffeas \add_in_i_a[6] (
	.clk(clk),
	.d(data_1_imag_i[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[6]~q ),
	.prn(vcc));
defparam \add_in_i_a[6] .is_wysiwyg = "true";
defparam \add_in_i_a[6] .power_up = "low";

dffeas \add_in_r_b[7] (
	.clk(clk),
	.d(data_3_real_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[7]~q ),
	.prn(vcc));
defparam \add_in_r_b[7] .is_wysiwyg = "true";
defparam \add_in_r_b[7] .power_up = "low";

dffeas \add_in_r_a[7] (
	.clk(clk),
	.d(data_1_real_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[7]~q ),
	.prn(vcc));
defparam \add_in_r_a[7] .is_wysiwyg = "true";
defparam \add_in_r_a[7] .power_up = "low";

dffeas \add_in_i_b[7] (
	.clk(clk),
	.d(data_3_imag_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[7]~q ),
	.prn(vcc));
defparam \add_in_i_b[7] .is_wysiwyg = "true";
defparam \add_in_i_b[7] .power_up = "low";

dffeas \add_in_i_a[7] (
	.clk(clk),
	.d(data_1_imag_i[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[7]~q ),
	.prn(vcc));
defparam \add_in_i_a[7] .is_wysiwyg = "true";
defparam \add_in_i_a[7] .power_up = "low";

dffeas \offset_counter[5] (
	.clk(clk),
	.d(\offset_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\offset_counter[5]~q ),
	.prn(vcc));
defparam \offset_counter[5] .is_wysiwyg = "true";
defparam \offset_counter[5] .power_up = "low";

dffeas \add_in_r_b[1] (
	.clk(clk),
	.d(data_3_real_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[1]~q ),
	.prn(vcc));
defparam \add_in_r_b[1] .is_wysiwyg = "true";
defparam \add_in_r_b[1] .power_up = "low";

dffeas \add_in_r_a[1] (
	.clk(clk),
	.d(data_1_real_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[1]~q ),
	.prn(vcc));
defparam \add_in_r_a[1] .is_wysiwyg = "true";
defparam \add_in_r_a[1] .power_up = "low";

dffeas \offset_counter[4] (
	.clk(clk),
	.d(\offset_counter~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\offset_counter[4]~q ),
	.prn(vcc));
defparam \offset_counter[4] .is_wysiwyg = "true";
defparam \offset_counter[4] .power_up = "low";

dffeas \add_in_i_b[1] (
	.clk(clk),
	.d(data_3_imag_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[1]~q ),
	.prn(vcc));
defparam \add_in_i_b[1] .is_wysiwyg = "true";
defparam \add_in_i_b[1] .power_up = "low";

dffeas \add_in_i_a[1] (
	.clk(clk),
	.d(data_1_imag_i[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[1]~q ),
	.prn(vcc));
defparam \add_in_i_a[1] .is_wysiwyg = "true";
defparam \add_in_i_a[1] .power_up = "low";

dffeas \offset_counter[3] (
	.clk(clk),
	.d(\offset_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\offset_counter[3]~q ),
	.prn(vcc));
defparam \offset_counter[3] .is_wysiwyg = "true";
defparam \offset_counter[3] .power_up = "low";

dffeas \offset_counter[2] (
	.clk(clk),
	.d(\offset_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\offset_counter[2]~q ),
	.prn(vcc));
defparam \offset_counter[2] .is_wysiwyg = "true";
defparam \offset_counter[2] .power_up = "low";

dffeas \offset_counter[0] (
	.clk(clk),
	.d(\offset_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\offset_counter[0]~q ),
	.prn(vcc));
defparam \offset_counter[0] .is_wysiwyg = "true";
defparam \offset_counter[0] .power_up = "low";

dffeas \offset_counter[1] (
	.clk(clk),
	.d(\offset_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\offset_counter[1]~q ),
	.prn(vcc));
defparam \offset_counter[1] .is_wysiwyg = "true";
defparam \offset_counter[1] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\offset_counter[3]~q ),
	.datab(!\offset_counter[2]~q ),
	.datac(!\offset_counter[0]~q ),
	.datad(!\offset_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \offset_counter~0 (
	.dataa(!reset_n),
	.datab(!tdl_arr_4),
	.datac(!\offset_counter[5]~q ),
	.datad(!\offset_counter[4]~q ),
	.datae(!\Add0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_counter~0 .extended_lut = "off";
defparam \offset_counter~0 .lut_mask = 64'hF77F7FF7F77F7FF7;
defparam \offset_counter~0 .shared_arith = "off";

dffeas \add_in_r_b[0] (
	.clk(clk),
	.d(data_3_real_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_b[0]~q ),
	.prn(vcc));
defparam \add_in_r_b[0] .is_wysiwyg = "true";
defparam \add_in_r_b[0] .power_up = "low";

dffeas \add_in_r_a[0] (
	.clk(clk),
	.d(data_1_real_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_r_a[0]~q ),
	.prn(vcc));
defparam \add_in_r_a[0] .is_wysiwyg = "true";
defparam \add_in_r_a[0] .power_up = "low";

cyclonev_lcell_comb \offset_counter~1 (
	.dataa(!reset_n),
	.datab(!tdl_arr_4),
	.datac(!\offset_counter[4]~q ),
	.datad(!\Add0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_counter~1 .extended_lut = "off";
defparam \offset_counter~1 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \offset_counter~1 .shared_arith = "off";

dffeas \add_in_i_b[0] (
	.clk(clk),
	.d(data_3_imag_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_b[0]~q ),
	.prn(vcc));
defparam \add_in_i_b[0] .is_wysiwyg = "true";
defparam \add_in_i_b[0] .power_up = "low";

dffeas \add_in_i_a[0] (
	.clk(clk),
	.d(data_1_imag_i[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\add_in_i_a[0]~q ),
	.prn(vcc));
defparam \add_in_i_a[0] .is_wysiwyg = "true";
defparam \add_in_i_a[0] .power_up = "low";

cyclonev_lcell_comb \offset_counter~2 (
	.dataa(!reset_n),
	.datab(!tdl_arr_4),
	.datac(!\offset_counter[3]~q ),
	.datad(!\offset_counter[2]~q ),
	.datae(!\offset_counter[0]~q ),
	.dataf(!\offset_counter[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_counter~2 .extended_lut = "off";
defparam \offset_counter~2 .lut_mask = 64'h7FF7F77FF77F7FF7;
defparam \offset_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \offset_counter~3 (
	.dataa(!reset_n),
	.datab(!tdl_arr_4),
	.datac(!\offset_counter[2]~q ),
	.datad(!\offset_counter[0]~q ),
	.datae(!\offset_counter[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_counter~3 .extended_lut = "off";
defparam \offset_counter~3 .lut_mask = 64'hF77F7FF7F77F7FF7;
defparam \offset_counter~3 .shared_arith = "off";

cyclonev_lcell_comb \offset_counter~4 (
	.dataa(!reset_n),
	.datab(!tdl_arr_4),
	.datac(!\offset_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_counter~4 .extended_lut = "off";
defparam \offset_counter~4 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \offset_counter~4 .shared_arith = "off";

cyclonev_lcell_comb \offset_counter~5 (
	.dataa(!reset_n),
	.datab(!tdl_arr_4),
	.datac(!\offset_counter[0]~q ),
	.datad(!\offset_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\offset_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \offset_counter~5 .extended_lut = "off";
defparam \offset_counter~5 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \offset_counter~5 .shared_arith = "off";

cyclonev_lcell_comb \sign_vec[1]~0 (
	.dataa(!\sign_sel[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sign_vec[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sign_vec[1]~0 .extended_lut = "off";
defparam \sign_vec[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sign_vec[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \sign_vec[3]~2 (
	.dataa(!\sign_sel[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sign_vec[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sign_vec[3]~2 .extended_lut = "off";
defparam \sign_vec[3]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sign_vec[3]~2 .shared_arith = "off";

dffeas \data_real_o[0] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_0),
	.prn(vcc));
defparam \data_real_o[0] .is_wysiwyg = "true";
defparam \data_real_o[0] .power_up = "low";

dffeas \data_real_o[1] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_1),
	.prn(vcc));
defparam \data_real_o[1] .is_wysiwyg = "true";
defparam \data_real_o[1] .power_up = "low";

dffeas \data_real_o[2] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_2),
	.prn(vcc));
defparam \data_real_o[2] .is_wysiwyg = "true";
defparam \data_real_o[2] .power_up = "low";

dffeas \data_real_o[3] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_3),
	.prn(vcc));
defparam \data_real_o[3] .is_wysiwyg = "true";
defparam \data_real_o[3] .power_up = "low";

dffeas \data_real_o[4] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_4),
	.prn(vcc));
defparam \data_real_o[4] .is_wysiwyg = "true";
defparam \data_real_o[4] .power_up = "low";

dffeas \data_real_o[5] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_5),
	.prn(vcc));
defparam \data_real_o[5] .is_wysiwyg = "true";
defparam \data_real_o[5] .power_up = "low";

dffeas \data_real_o[6] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_6),
	.prn(vcc));
defparam \data_real_o[6] .is_wysiwyg = "true";
defparam \data_real_o[6] .power_up = "low";

dffeas \data_real_o[7] (
	.clk(clk),
	.d(\gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(data_real_o_7),
	.prn(vcc));
defparam \data_real_o[7] .is_wysiwyg = "true";
defparam \data_real_o[7] .power_up = "low";

dffeas \data_imag_o[0] (
	.clk(clk),
	.d(\data_imag_o[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_0),
	.prn(vcc));
defparam \data_imag_o[0] .is_wysiwyg = "true";
defparam \data_imag_o[0] .power_up = "low";

dffeas \data_imag_o[1] (
	.clk(clk),
	.d(\data_imag_o[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_1),
	.prn(vcc));
defparam \data_imag_o[1] .is_wysiwyg = "true";
defparam \data_imag_o[1] .power_up = "low";

dffeas \data_imag_o[2] (
	.clk(clk),
	.d(\data_imag_o[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_2),
	.prn(vcc));
defparam \data_imag_o[2] .is_wysiwyg = "true";
defparam \data_imag_o[2] .power_up = "low";

dffeas \data_imag_o[3] (
	.clk(clk),
	.d(\data_imag_o[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_3),
	.prn(vcc));
defparam \data_imag_o[3] .is_wysiwyg = "true";
defparam \data_imag_o[3] .power_up = "low";

dffeas \data_imag_o[4] (
	.clk(clk),
	.d(\data_imag_o[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_4),
	.prn(vcc));
defparam \data_imag_o[4] .is_wysiwyg = "true";
defparam \data_imag_o[4] .power_up = "low";

dffeas \data_imag_o[5] (
	.clk(clk),
	.d(\data_imag_o[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_5),
	.prn(vcc));
defparam \data_imag_o[5] .is_wysiwyg = "true";
defparam \data_imag_o[5] .power_up = "low";

dffeas \data_imag_o[6] (
	.clk(clk),
	.d(\data_imag_o[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_6),
	.prn(vcc));
defparam \data_imag_o[6] .is_wysiwyg = "true";
defparam \data_imag_o[6] .power_up = "low";

dffeas \data_imag_o[7] (
	.clk(clk),
	.d(\data_imag_o[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_imag_o_7),
	.prn(vcc));
defparam \data_imag_o[7] .is_wysiwyg = "true";
defparam \data_imag_o[7] .power_up = "low";

cyclonev_lcell_comb \data_imag_o[0]~0 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_0),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[0]~0 .extended_lut = "off";
defparam \data_imag_o[0]~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[1]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_1),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[1]~1 .extended_lut = "off";
defparam \data_imag_o[1]~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[2]~2 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_2),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[2]~2 .extended_lut = "off";
defparam \data_imag_o[2]~2 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[3]~3 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_3),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[3]~3 .extended_lut = "off";
defparam \data_imag_o[3]~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[4]~4 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_4),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[4]~4 .extended_lut = "off";
defparam \data_imag_o[4]~4 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[5]~5 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_5),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[5]~5 .extended_lut = "off";
defparam \data_imag_o[5]~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[6]~6 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_6),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[6]~6 .extended_lut = "off";
defparam \data_imag_o[6]~6 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \data_imag_o[7]~7 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!data_imag_o_7),
	.datad(!\gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_imag_o[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_imag_o[7]~7 .extended_lut = "off";
defparam \data_imag_o[7]~7 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \data_imag_o[7]~7 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_14 (
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	output_r_2,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	output_r_8,
	output_r_9,
	output_r_1,
	output_r_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	output_r_2;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	output_r_8;
input 	output_r_9;
input 	output_r_1;
input 	output_r_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_15 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.output_r_2(output_r_2),
	.output_r_3(output_r_3),
	.output_r_4(output_r_4),
	.output_r_5(output_r_5),
	.output_r_6(output_r_6),
	.output_r_7(output_r_7),
	.output_r_8(output_r_8),
	.output_r_9(output_r_9),
	.output_r_1(output_r_1),
	.output_r_0(output_r_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_15 (
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	output_r_2,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	output_r_8,
	output_r_9,
	output_r_1,
	output_r_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	output_r_2;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	output_r_8;
input 	output_r_9;
input 	output_r_1;
input 	output_r_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_8 auto_generated(
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.output_r_2(output_r_2),
	.output_r_3(output_r_3),
	.output_r_4(output_r_4),
	.output_r_5(output_r_5),
	.output_r_6(output_r_6),
	.output_r_7(output_r_7),
	.output_r_8(output_r_8),
	.output_r_9(output_r_9),
	.output_r_1(output_r_1),
	.output_r_0(output_r_0),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_8 (
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	output_r_2,
	output_r_3,
	output_r_4,
	output_r_5,
	output_r_6,
	output_r_7,
	output_r_8,
	output_r_9,
	output_r_1,
	output_r_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	output_r_2;
input 	output_r_3;
input 	output_r_4;
input 	output_r_5;
input 	output_r_6;
input 	output_r_7;
input 	output_r_8;
input 	output_r_9;
input 	output_r_1;
input 	output_r_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_r_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u0|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_pround_15 (
	global_clock_enable,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	output_i_2,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	output_i_8,
	output_i_9,
	output_i_1,
	output_i_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	output_i_2;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	output_i_8;
input 	output_i_9;
input 	output_i_1;
input 	output_i_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_LPM_ADD_SUB_16 \gbrnd:nev:gp:lpm_add_sub_component (
	.clken(global_clock_enable),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.output_i_2(output_i_2),
	.output_i_3(output_i_3),
	.output_i_4(output_i_4),
	.output_i_5(output_i_5),
	.output_i_6(output_i_6),
	.output_i_7(output_i_7),
	.output_i_8(output_i_8),
	.output_i_9(output_i_9),
	.output_i_1(output_i_1),
	.output_i_0(output_i_0),
	.clock(clk));

endmodule

module IFFT_LPM_ADD_SUB_16 (
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	output_i_2,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	output_i_8,
	output_i_9,
	output_i_1,
	output_i_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	output_i_2;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	output_i_8;
input 	output_i_9;
input 	output_i_1;
input 	output_i_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_add_sub_2gj_9 auto_generated(
	.clken(clken),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.output_i_2(output_i_2),
	.output_i_3(output_i_3),
	.output_i_4(output_i_4),
	.output_i_5(output_i_5),
	.output_i_6(output_i_6),
	.output_i_7(output_i_7),
	.output_i_8(output_i_8),
	.output_i_9(output_i_9),
	.output_i_1(output_i_1),
	.output_i_0(output_i_0),
	.clock(clock));

endmodule

module IFFT_add_sub_2gj_9 (
	clken,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	output_i_2,
	output_i_3,
	output_i_4,
	output_i_5,
	output_i_6,
	output_i_7,
	output_i_8,
	output_i_9,
	output_i_1,
	output_i_0,
	clock)/* synthesis synthesis_greybox=1 */;
input 	clken;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	output_i_2;
input 	output_i_3;
input 	output_i_4;
input 	output_i_5;
input 	output_i_6;
input 	output_i_7;
input 	output_i_8;
input 	output_i_9;
input 	output_i_1;
input 	output_i_0;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ;
wire \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ;


dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .lut_mask = 64'h000000000000FF00;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25_sumout ),
	.cout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!output_i_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29_sumout ),
	.cout(),
	.shareout());
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .extended_lut = "off";
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .lut_mask = 64'h00000000000000FF;
defparam \fft_ii_0|asj_fft_sglstream_inst|gen_radix_4_last_pass:lpp|gen_full_rnd:u1|gbrnd:nev:gp:lpm_add_sub_component|auto_generated|op_1~29 .shared_arith = "off";

endmodule

module IFFT_asj_fft_lpprdadgen (
	tdl_arr_4,
	tdl_arr_19,
	data_rdy_int,
	tdl_arr_0_4,
	tdl_arr_1_4,
	global_clock_enable,
	rd_addr_d_0,
	rd_addr_d_1,
	sw_0,
	sw_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_4;
input 	tdl_arr_19;
input 	data_rdy_int;
output 	tdl_arr_0_4;
output 	tdl_arr_1_4;
input 	global_clock_enable;
output 	rd_addr_d_0;
output 	rd_addr_d_1;
output 	sw_0;
output 	sw_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \en_d~q ;
wire \en_i~0_combout ;
wire \en_i~q ;
wire \count~2_combout ;
wire \count[0]~q ;
wire \count~3_combout ;
wire \count[1]~q ;
wire \count~0_combout ;
wire \count[2]~q ;
wire \count~1_combout ;
wire \count[3]~q ;
wire \Add1~0_combout ;
wire \Add1~1_combout ;


IFFT_asj_fft_tdl_rst \gen_M4K:delay_swd (
	.tdl_arr_0_4(tdl_arr_0_4),
	.tdl_arr_1_4(tdl_arr_1_4),
	.global_clock_enable(global_clock_enable),
	.sw_0(sw_0),
	.sw_1(sw_1),
	.clk(clk),
	.reset_n(reset_n));

IFFT_asj_fft_tdl_bit_rst_4 delay_en(
	.tdl_arr_4(tdl_arr_4),
	.en_i(\en_i~q ),
	.global_clock_enable(global_clock_enable),
	.clk(clk),
	.reset_n(reset_n));

dffeas \rd_addr_d[0] (
	.clk(clk),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_d_0),
	.prn(vcc));
defparam \rd_addr_d[0] .is_wysiwyg = "true";
defparam \rd_addr_d[0] .power_up = "low";

dffeas \rd_addr_d[1] (
	.clk(clk),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(rd_addr_d_1),
	.prn(vcc));
defparam \rd_addr_d[1] .is_wysiwyg = "true";
defparam \rd_addr_d[1] .power_up = "low";

dffeas \sw[0] (
	.clk(clk),
	.d(\Add1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(sw_0),
	.prn(vcc));
defparam \sw[0] .is_wysiwyg = "true";
defparam \sw[0] .power_up = "low";

dffeas \sw[1] (
	.clk(clk),
	.d(\Add1~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(sw_1),
	.prn(vcc));
defparam \sw[1] .is_wysiwyg = "true";
defparam \sw[1] .power_up = "low";

dffeas en_d(
	.clk(clk),
	.d(tdl_arr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\en_d~q ),
	.prn(vcc));
defparam en_d.is_wysiwyg = "true";
defparam en_d.power_up = "low";

cyclonev_lcell_comb \en_i~0 (
	.dataa(!\en_d~q ),
	.datab(!tdl_arr_19),
	.datac(!data_rdy_int),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\en_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \en_i~0 .extended_lut = "off";
defparam \en_i~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \en_i~0 .shared_arith = "off";

dffeas en_i(
	.clk(clk),
	.d(\en_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\en_i~q ),
	.prn(vcc));
defparam en_i.is_wysiwyg = "true";
defparam en_i.power_up = "low";

cyclonev_lcell_comb \count~2 (
	.dataa(!reset_n),
	.datab(!\en_i~q ),
	.datac(!\count[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~2 .extended_lut = "off";
defparam \count~2 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \count~2 .shared_arith = "off";

dffeas \count[0] (
	.clk(clk),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclonev_lcell_comb \count~3 (
	.dataa(!reset_n),
	.datab(!\en_i~q ),
	.datac(!\count[0]~q ),
	.datad(!\count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~3 .extended_lut = "off";
defparam \count~3 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \count~3 .shared_arith = "off";

dffeas \count[1] (
	.clk(clk),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \count~0 (
	.dataa(!reset_n),
	.datab(!\en_i~q ),
	.datac(!\count[2]~q ),
	.datad(!\count[0]~q ),
	.datae(!\count[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~0 .extended_lut = "off";
defparam \count~0 .lut_mask = 64'hFDDFDFFDFDDFDFFD;
defparam \count~0 .shared_arith = "off";

dffeas \count[2] (
	.clk(clk),
	.d(\count~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cyclonev_lcell_comb \count~1 (
	.dataa(!reset_n),
	.datab(!\en_i~q ),
	.datac(!\count[2]~q ),
	.datad(!\count[3]~q ),
	.datae(!\count[0]~q ),
	.dataf(!\count[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~1 .extended_lut = "off";
defparam \count~1 .lut_mask = 64'hDFFDFDDFFDDFDFFD;
defparam \count~1 .shared_arith = "off";

dffeas \count[3] (
	.clk(clk),
	.d(\count~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\count[2]~q ),
	.datab(!\count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h6666666666666666;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\count[2]~q ),
	.datab(!\count[3]~q ),
	.datac(!\count[0]~q ),
	.datad(!\count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h6996699669966996;
defparam \Add1~1 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl_bit_rst_4 (
	tdl_arr_4,
	en_i,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_4;
input 	en_i;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;


dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_4),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(en_i),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_rst (
	tdl_arr_0_4,
	tdl_arr_1_4,
	global_clock_enable,
	sw_0,
	sw_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_0_4;
output 	tdl_arr_1_4;
input 	global_clock_enable;
input 	sw_0;
input 	sw_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0][0]~q ;
wire \tdl_arr[1][0]~q ;
wire \tdl_arr[2][0]~q ;
wire \tdl_arr[3][0]~q ;
wire \tdl_arr[0][1]~q ;
wire \tdl_arr[1][1]~q ;
wire \tdl_arr[2][1]~q ;
wire \tdl_arr[3][1]~q ;


dffeas \tdl_arr[4][0] (
	.clk(clk),
	.d(\tdl_arr[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_0_4),
	.prn(vcc));
defparam \tdl_arr[4][0] .is_wysiwyg = "true";
defparam \tdl_arr[4][0] .power_up = "low";

dffeas \tdl_arr[4][1] (
	.clk(clk),
	.d(\tdl_arr[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_1_4),
	.prn(vcc));
defparam \tdl_arr[4][1] .is_wysiwyg = "true";
defparam \tdl_arr[4][1] .power_up = "low";

dffeas \tdl_arr[0][0] (
	.clk(clk),
	.d(sw_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][0]~q ),
	.prn(vcc));
defparam \tdl_arr[0][0] .is_wysiwyg = "true";
defparam \tdl_arr[0][0] .power_up = "low";

dffeas \tdl_arr[1][0] (
	.clk(clk),
	.d(\tdl_arr[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1][0]~q ),
	.prn(vcc));
defparam \tdl_arr[1][0] .is_wysiwyg = "true";
defparam \tdl_arr[1][0] .power_up = "low";

dffeas \tdl_arr[2][0] (
	.clk(clk),
	.d(\tdl_arr[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2][0]~q ),
	.prn(vcc));
defparam \tdl_arr[2][0] .is_wysiwyg = "true";
defparam \tdl_arr[2][0] .power_up = "low";

dffeas \tdl_arr[3][0] (
	.clk(clk),
	.d(\tdl_arr[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3][0]~q ),
	.prn(vcc));
defparam \tdl_arr[3][0] .is_wysiwyg = "true";
defparam \tdl_arr[3][0] .power_up = "low";

dffeas \tdl_arr[0][1] (
	.clk(clk),
	.d(sw_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0][1]~q ),
	.prn(vcc));
defparam \tdl_arr[0][1] .is_wysiwyg = "true";
defparam \tdl_arr[0][1] .power_up = "low";

dffeas \tdl_arr[1][1] (
	.clk(clk),
	.d(\tdl_arr[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1][1]~q ),
	.prn(vcc));
defparam \tdl_arr[1][1] .is_wysiwyg = "true";
defparam \tdl_arr[1][1] .power_up = "low";

dffeas \tdl_arr[2][1] (
	.clk(clk),
	.d(\tdl_arr[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2][1]~q ),
	.prn(vcc));
defparam \tdl_arr[2][1] .is_wysiwyg = "true";
defparam \tdl_arr[2][1] .power_up = "low";

dffeas \tdl_arr[3][1] (
	.clk(clk),
	.d(\tdl_arr[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3][1]~q ),
	.prn(vcc));
defparam \tdl_arr[3][1] .is_wysiwyg = "true";
defparam \tdl_arr[3][1] .power_up = "low";

endmodule

module IFFT_asj_fft_m_k_counter (
	blk_done_int1,
	next_block,
	p_0,
	data_rdy_vec_4,
	next_pass_i1,
	global_clock_enable,
	p_1,
	k_count_1,
	k_count_3,
	k_count_0,
	k_count_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	blk_done_int1;
input 	next_block;
output 	p_0;
input 	data_rdy_vec_4;
output 	next_pass_i1;
input 	global_clock_enable;
output 	p_1;
output 	k_count_1;
output 	k_count_3;
output 	k_count_0;
output 	k_count_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \next_block_d~q ;
wire \next_block_d2~q ;
wire \next_block_d3~q ;
wire \next_block_d4~q ;
wire \k_state.HOLD~0_combout ;
wire \k_state.HOLD~q ;
wire \del_npi_cnt~1_combout ;
wire \del_npi_cnt[0]~q ;
wire \del_npi_cnt~2_combout ;
wire \del_npi_cnt[1]~q ;
wire \del_npi_cnt~3_combout ;
wire \del_npi_cnt[2]~q ;
wire \del_npi_cnt~4_combout ;
wire \del_npi_cnt[3]~q ;
wire \del_npi_cnt~5_combout ;
wire \del_npi_cnt[4]~q ;
wire \next_pass_id~0_combout ;
wire \next_pass_id~1_combout ;
wire \next_pass_id~q ;
wire \k~0_combout ;
wire \k_state~8_combout ;
wire \k_state.IDLE~q ;
wire \k[0]~1_combout ;
wire \k[0]~q ;
wire \k~2_combout ;
wire \k[1]~q ;
wire \k~3_combout ;
wire \k[2]~q ;
wire \k~4_combout ;
wire \k[3]~q ;
wire \k_state~7_combout ;
wire \Selector0~0_combout ;
wire \k_state.RUN_CNT~q ;
wire \k_state~6_combout ;
wire \k_state.NEXT_PASS_UPD~q ;
wire \blk_done_int~0_combout ;
wire \p~2_combout ;
wire \p[0]~1_combout ;
wire \p~0_combout ;


dffeas blk_done_int(
	.clk(clk),
	.d(\blk_done_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(blk_done_int1),
	.prn(vcc));
defparam blk_done_int.is_wysiwyg = "true";
defparam blk_done_int.power_up = "low";

dffeas \p[0] (
	.clk(clk),
	.d(\p~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\p[0]~1_combout ),
	.q(p_0),
	.prn(vcc));
defparam \p[0] .is_wysiwyg = "true";
defparam \p[0] .power_up = "low";

dffeas next_pass_i(
	.clk(clk),
	.d(\k_state.NEXT_PASS_UPD~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(next_pass_i1),
	.prn(vcc));
defparam next_pass_i.is_wysiwyg = "true";
defparam next_pass_i.power_up = "low";

dffeas \p[1] (
	.clk(clk),
	.d(\p~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\p[0]~1_combout ),
	.q(p_1),
	.prn(vcc));
defparam \p[1] .is_wysiwyg = "true";
defparam \p[1] .power_up = "low";

dffeas \k_count[1] (
	.clk(clk),
	.d(\k[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(k_count_1),
	.prn(vcc));
defparam \k_count[1] .is_wysiwyg = "true";
defparam \k_count[1] .power_up = "low";

dffeas \k_count[3] (
	.clk(clk),
	.d(\k[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(k_count_3),
	.prn(vcc));
defparam \k_count[3] .is_wysiwyg = "true";
defparam \k_count[3] .power_up = "low";

dffeas \k_count[0] (
	.clk(clk),
	.d(\k[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(k_count_0),
	.prn(vcc));
defparam \k_count[0] .is_wysiwyg = "true";
defparam \k_count[0] .power_up = "low";

dffeas \k_count[2] (
	.clk(clk),
	.d(\k[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(k_count_2),
	.prn(vcc));
defparam \k_count[2] .is_wysiwyg = "true";
defparam \k_count[2] .power_up = "low";

dffeas next_block_d(
	.clk(clk),
	.d(next_block),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\next_block_d~q ),
	.prn(vcc));
defparam next_block_d.is_wysiwyg = "true";
defparam next_block_d.power_up = "low";

dffeas next_block_d2(
	.clk(clk),
	.d(\next_block_d~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\next_block_d2~q ),
	.prn(vcc));
defparam next_block_d2.is_wysiwyg = "true";
defparam next_block_d2.power_up = "low";

dffeas next_block_d3(
	.clk(clk),
	.d(\next_block_d2~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\next_block_d3~q ),
	.prn(vcc));
defparam next_block_d3.is_wysiwyg = "true";
defparam next_block_d3.power_up = "low";

dffeas next_block_d4(
	.clk(clk),
	.d(\next_block_d3~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\next_block_d4~q ),
	.prn(vcc));
defparam next_block_d4.is_wysiwyg = "true";
defparam next_block_d4.power_up = "low";

cyclonev_lcell_comb \k_state.HOLD~0 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\k_state.NEXT_PASS_UPD~q ),
	.datad(!\next_block_d4~q ),
	.datae(!\next_pass_id~q ),
	.dataf(!\k_state.HOLD~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k_state.HOLD~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k_state.HOLD~0 .extended_lut = "off";
defparam \k_state.HOLD~0 .lut_mask = 64'hFF7FDF5FFFFFFFFF;
defparam \k_state.HOLD~0 .shared_arith = "off";

dffeas \k_state.HOLD (
	.clk(clk),
	.d(\k_state.HOLD~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\k_state.HOLD~q ),
	.prn(vcc));
defparam \k_state.HOLD .is_wysiwyg = "true";
defparam \k_state.HOLD .power_up = "low";

cyclonev_lcell_comb \del_npi_cnt~1 (
	.dataa(!\k_state.HOLD~q ),
	.datab(!\del_npi_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_npi_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_npi_cnt~1 .extended_lut = "off";
defparam \del_npi_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \del_npi_cnt~1 .shared_arith = "off";

dffeas \del_npi_cnt[0] (
	.clk(clk),
	.d(\del_npi_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_npi_cnt[0]~q ),
	.prn(vcc));
defparam \del_npi_cnt[0] .is_wysiwyg = "true";
defparam \del_npi_cnt[0] .power_up = "low";

cyclonev_lcell_comb \del_npi_cnt~2 (
	.dataa(!\k_state.HOLD~q ),
	.datab(!\del_npi_cnt[0]~q ),
	.datac(!\del_npi_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_npi_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_npi_cnt~2 .extended_lut = "off";
defparam \del_npi_cnt~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \del_npi_cnt~2 .shared_arith = "off";

dffeas \del_npi_cnt[1] (
	.clk(clk),
	.d(\del_npi_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_npi_cnt[1]~q ),
	.prn(vcc));
defparam \del_npi_cnt[1] .is_wysiwyg = "true";
defparam \del_npi_cnt[1] .power_up = "low";

cyclonev_lcell_comb \del_npi_cnt~3 (
	.dataa(!\k_state.HOLD~q ),
	.datab(!\del_npi_cnt[2]~q ),
	.datac(!\del_npi_cnt[0]~q ),
	.datad(!\del_npi_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_npi_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_npi_cnt~3 .extended_lut = "off";
defparam \del_npi_cnt~3 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \del_npi_cnt~3 .shared_arith = "off";

dffeas \del_npi_cnt[2] (
	.clk(clk),
	.d(\del_npi_cnt~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_npi_cnt[2]~q ),
	.prn(vcc));
defparam \del_npi_cnt[2] .is_wysiwyg = "true";
defparam \del_npi_cnt[2] .power_up = "low";

cyclonev_lcell_comb \del_npi_cnt~4 (
	.dataa(!\k_state.HOLD~q ),
	.datab(!\del_npi_cnt[2]~q ),
	.datac(!\del_npi_cnt[3]~q ),
	.datad(!\del_npi_cnt[0]~q ),
	.datae(!\del_npi_cnt[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_npi_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_npi_cnt~4 .extended_lut = "off";
defparam \del_npi_cnt~4 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \del_npi_cnt~4 .shared_arith = "off";

dffeas \del_npi_cnt[3] (
	.clk(clk),
	.d(\del_npi_cnt~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_npi_cnt[3]~q ),
	.prn(vcc));
defparam \del_npi_cnt[3] .is_wysiwyg = "true";
defparam \del_npi_cnt[3] .power_up = "low";

cyclonev_lcell_comb \del_npi_cnt~5 (
	.dataa(!\k_state.HOLD~q ),
	.datab(!\del_npi_cnt[2]~q ),
	.datac(!\del_npi_cnt[3]~q ),
	.datad(!\del_npi_cnt[4]~q ),
	.datae(!\del_npi_cnt[0]~q ),
	.dataf(!\del_npi_cnt[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\del_npi_cnt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \del_npi_cnt~5 .extended_lut = "off";
defparam \del_npi_cnt~5 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \del_npi_cnt~5 .shared_arith = "off";

dffeas \del_npi_cnt[4] (
	.clk(clk),
	.d(\del_npi_cnt~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\del_npi_cnt[4]~q ),
	.prn(vcc));
defparam \del_npi_cnt[4] .is_wysiwyg = "true";
defparam \del_npi_cnt[4] .power_up = "low";

cyclonev_lcell_comb \next_pass_id~0 (
	.dataa(!\k_state.HOLD~q ),
	.datab(!\del_npi_cnt[2]~q ),
	.datac(!\del_npi_cnt[3]~q ),
	.datad(!\del_npi_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\next_pass_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \next_pass_id~0 .extended_lut = "off";
defparam \next_pass_id~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \next_pass_id~0 .shared_arith = "off";

cyclonev_lcell_comb \next_pass_id~1 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!\del_npi_cnt[0]~q ),
	.datad(!\del_npi_cnt[1]~q ),
	.datae(!\next_pass_id~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\next_pass_id~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \next_pass_id~1 .extended_lut = "off";
defparam \next_pass_id~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \next_pass_id~1 .shared_arith = "off";

dffeas next_pass_id(
	.clk(clk),
	.d(\next_pass_id~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\next_pass_id~q ),
	.prn(vcc));
defparam next_pass_id.is_wysiwyg = "true";
defparam next_pass_id.power_up = "low";

cyclonev_lcell_comb \k~0 (
	.dataa(!reset_n),
	.datab(!next_block),
	.datac(!\k[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k~0 .extended_lut = "off";
defparam \k~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \k~0 .shared_arith = "off";

cyclonev_lcell_comb \k_state~8 (
	.dataa(!reset_n),
	.datab(!\next_block_d4~q ),
	.datac(!\k_state.IDLE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k_state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k_state~8 .extended_lut = "off";
defparam \k_state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \k_state~8 .shared_arith = "off";

dffeas \k_state.IDLE (
	.clk(clk),
	.d(\k_state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\k_state.IDLE~q ),
	.prn(vcc));
defparam \k_state.IDLE .is_wysiwyg = "true";
defparam \k_state.IDLE .power_up = "low";

cyclonev_lcell_comb \k[0]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!next_block),
	.datad(!\k_state.HOLD~q ),
	.datae(!\k_state.IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k[0]~1 .extended_lut = "off";
defparam \k[0]~1 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \k[0]~1 .shared_arith = "off";

dffeas \k[0] (
	.clk(clk),
	.d(\k~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\k[0]~1_combout ),
	.q(\k[0]~q ),
	.prn(vcc));
defparam \k[0] .is_wysiwyg = "true";
defparam \k[0] .power_up = "low";

cyclonev_lcell_comb \k~2 (
	.dataa(!reset_n),
	.datab(!next_block),
	.datac(!\k[0]~q ),
	.datad(!\k[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k~2 .extended_lut = "off";
defparam \k~2 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \k~2 .shared_arith = "off";

dffeas \k[1] (
	.clk(clk),
	.d(\k~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\k[0]~1_combout ),
	.q(\k[1]~q ),
	.prn(vcc));
defparam \k[1] .is_wysiwyg = "true";
defparam \k[1] .power_up = "low";

cyclonev_lcell_comb \k~3 (
	.dataa(!reset_n),
	.datab(!next_block),
	.datac(!\k[0]~q ),
	.datad(!\k[1]~q ),
	.datae(!\k[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k~3 .extended_lut = "off";
defparam \k~3 .lut_mask = 64'hFDDFDFFDFDDFDFFD;
defparam \k~3 .shared_arith = "off";

dffeas \k[2] (
	.clk(clk),
	.d(\k~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\k[0]~1_combout ),
	.q(\k[2]~q ),
	.prn(vcc));
defparam \k[2] .is_wysiwyg = "true";
defparam \k[2] .power_up = "low";

cyclonev_lcell_comb \k~4 (
	.dataa(!reset_n),
	.datab(!next_block),
	.datac(!\k[0]~q ),
	.datad(!\k[1]~q ),
	.datae(!\k[2]~q ),
	.dataf(!\k[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k~4 .extended_lut = "off";
defparam \k~4 .lut_mask = 64'hDFFDFDDFFDDFDFFD;
defparam \k~4 .shared_arith = "off";

dffeas \k[3] (
	.clk(clk),
	.d(\k~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\k[0]~1_combout ),
	.q(\k[3]~q ),
	.prn(vcc));
defparam \k[3] .is_wysiwyg = "true";
defparam \k[3] .power_up = "low";

cyclonev_lcell_comb \k_state~7 (
	.dataa(!\k[0]~q ),
	.datab(!\k[1]~q ),
	.datac(!\k[2]~q ),
	.datad(!\k[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k_state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k_state~7 .extended_lut = "off";
defparam \k_state~7 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \k_state~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\next_block_d4~q ),
	.datab(!\k_state.RUN_CNT~q ),
	.datac(!\next_pass_id~q ),
	.datad(!\k_state.HOLD~q ),
	.datae(!\k_state~7_combout ),
	.dataf(!\k_state.IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \Selector0~0 .shared_arith = "off";

dffeas \k_state.RUN_CNT (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\k_state.RUN_CNT~q ),
	.prn(vcc));
defparam \k_state.RUN_CNT .is_wysiwyg = "true";
defparam \k_state.RUN_CNT .power_up = "low";

cyclonev_lcell_comb \k_state~6 (
	.dataa(!reset_n),
	.datab(!\k_state.RUN_CNT~q ),
	.datac(!\k[0]~q ),
	.datad(!\k[1]~q ),
	.datae(!\k[2]~q ),
	.dataf(!\k[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\k_state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \k_state~6 .extended_lut = "off";
defparam \k_state~6 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \k_state~6 .shared_arith = "off";

dffeas \k_state.NEXT_PASS_UPD (
	.clk(clk),
	.d(\k_state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\k_state.NEXT_PASS_UPD~q ),
	.prn(vcc));
defparam \k_state.NEXT_PASS_UPD .is_wysiwyg = "true";
defparam \k_state.NEXT_PASS_UPD .power_up = "low";

cyclonev_lcell_comb \blk_done_int~0 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!\k_state.NEXT_PASS_UPD~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\blk_done_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \blk_done_int~0 .extended_lut = "off";
defparam \blk_done_int~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \blk_done_int~0 .shared_arith = "off";

cyclonev_lcell_comb \p~2 (
	.dataa(!p_1),
	.datab(!p_0),
	.datac(!\next_block_d4~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p~2 .extended_lut = "off";
defparam \p~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \p~2 .shared_arith = "off";

cyclonev_lcell_comb \p[0]~1 (
	.dataa(!reset_n),
	.datab(!global_clock_enable),
	.datac(!\next_block_d4~q ),
	.datad(!data_rdy_vec_4),
	.datae(!next_pass_i1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p[0]~1 .extended_lut = "off";
defparam \p[0]~1 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \p[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \p~0 (
	.dataa(!reset_n),
	.datab(!p_1),
	.datac(!p_0),
	.datad(!\next_block_d4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\p~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \p~0 .extended_lut = "off";
defparam \p~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \p~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_tdl_bit_rst_5 (
	blk_done_int,
	tdl_arr_11,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	blk_done_int;
output 	tdl_arr_11;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;
wire \tdl_arr[8]~q ;
wire \tdl_arr[9]~q ;
wire \tdl_arr[10]~q ;


dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_11),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(blk_done_int),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_bit_rst_6 (
	tdl_arr_11,
	tdl_arr_19,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	tdl_arr_11;
output 	tdl_arr_19;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;
wire \tdl_arr[8]~q ;
wire \tdl_arr[9]~q ;
wire \tdl_arr[10]~q ;
wire \tdl_arr[11]~q ;
wire \tdl_arr[12]~q ;
wire \tdl_arr[13]~q ;
wire \tdl_arr[14]~q ;
wire \tdl_arr[15]~q ;
wire \tdl_arr[16]~q ;
wire \tdl_arr[17]~q ;
wire \tdl_arr[18]~q ;


dffeas \tdl_arr[19] (
	.clk(clk),
	.d(\tdl_arr[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_19),
	.prn(vcc));
defparam \tdl_arr[19] .is_wysiwyg = "true";
defparam \tdl_arr[19] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(tdl_arr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[9]~q ),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[10] (
	.clk(clk),
	.d(\tdl_arr[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[10]~q ),
	.prn(vcc));
defparam \tdl_arr[10] .is_wysiwyg = "true";
defparam \tdl_arr[10] .power_up = "low";

dffeas \tdl_arr[11] (
	.clk(clk),
	.d(\tdl_arr[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[11]~q ),
	.prn(vcc));
defparam \tdl_arr[11] .is_wysiwyg = "true";
defparam \tdl_arr[11] .power_up = "low";

dffeas \tdl_arr[12] (
	.clk(clk),
	.d(\tdl_arr[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[12]~q ),
	.prn(vcc));
defparam \tdl_arr[12] .is_wysiwyg = "true";
defparam \tdl_arr[12] .power_up = "low";

dffeas \tdl_arr[13] (
	.clk(clk),
	.d(\tdl_arr[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[13]~q ),
	.prn(vcc));
defparam \tdl_arr[13] .is_wysiwyg = "true";
defparam \tdl_arr[13] .power_up = "low";

dffeas \tdl_arr[14] (
	.clk(clk),
	.d(\tdl_arr[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[14]~q ),
	.prn(vcc));
defparam \tdl_arr[14] .is_wysiwyg = "true";
defparam \tdl_arr[14] .power_up = "low";

dffeas \tdl_arr[15] (
	.clk(clk),
	.d(\tdl_arr[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[15]~q ),
	.prn(vcc));
defparam \tdl_arr[15] .is_wysiwyg = "true";
defparam \tdl_arr[15] .power_up = "low";

dffeas \tdl_arr[16] (
	.clk(clk),
	.d(\tdl_arr[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[16]~q ),
	.prn(vcc));
defparam \tdl_arr[16] .is_wysiwyg = "true";
defparam \tdl_arr[16] .power_up = "low";

dffeas \tdl_arr[17] (
	.clk(clk),
	.d(\tdl_arr[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[17]~q ),
	.prn(vcc));
defparam \tdl_arr[17] .is_wysiwyg = "true";
defparam \tdl_arr[17] .power_up = "low";

dffeas \tdl_arr[18] (
	.clk(clk),
	.d(\tdl_arr[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[18]~q ),
	.prn(vcc));
defparam \tdl_arr[18] .is_wysiwyg = "true";
defparam \tdl_arr[18] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_bit_rst_8 (
	next_pass_i,
	tdl_arr_9,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	next_pass_i;
output 	tdl_arr_9;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;
wire \tdl_arr[5]~q ;
wire \tdl_arr[6]~q ;
wire \tdl_arr[7]~q ;
wire \tdl_arr[8]~q ;


dffeas \tdl_arr[9] (
	.clk(clk),
	.d(\tdl_arr[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_9),
	.prn(vcc));
defparam \tdl_arr[9] .is_wysiwyg = "true";
defparam \tdl_arr[9] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(next_pass_i),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[5]~q ),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[6] (
	.clk(clk),
	.d(\tdl_arr[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[6]~q ),
	.prn(vcc));
defparam \tdl_arr[6] .is_wysiwyg = "true";
defparam \tdl_arr[6] .power_up = "low";

dffeas \tdl_arr[7] (
	.clk(clk),
	.d(\tdl_arr[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[7]~q ),
	.prn(vcc));
defparam \tdl_arr[7] .is_wysiwyg = "true";
defparam \tdl_arr[7] .power_up = "low";

dffeas \tdl_arr[8] (
	.clk(clk),
	.d(\tdl_arr[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[8]~q ),
	.prn(vcc));
defparam \tdl_arr[8] .is_wysiwyg = "true";
defparam \tdl_arr[8] .power_up = "low";

endmodule

module IFFT_asj_fft_tdl_bit_rst_9 (
	tdl_arr_5,
	tdl_arr_4,
	global_clock_enable,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdl_arr_5;
input 	tdl_arr_4;
input 	global_clock_enable;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \tdl_arr[0]~q ;
wire \tdl_arr[1]~q ;
wire \tdl_arr[2]~q ;
wire \tdl_arr[3]~q ;
wire \tdl_arr[4]~q ;


dffeas \tdl_arr[5] (
	.clk(clk),
	.d(\tdl_arr[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(tdl_arr_5),
	.prn(vcc));
defparam \tdl_arr[5] .is_wysiwyg = "true";
defparam \tdl_arr[5] .power_up = "low";

dffeas \tdl_arr[0] (
	.clk(clk),
	.d(tdl_arr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[0]~q ),
	.prn(vcc));
defparam \tdl_arr[0] .is_wysiwyg = "true";
defparam \tdl_arr[0] .power_up = "low";

dffeas \tdl_arr[1] (
	.clk(clk),
	.d(\tdl_arr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[1]~q ),
	.prn(vcc));
defparam \tdl_arr[1] .is_wysiwyg = "true";
defparam \tdl_arr[1] .power_up = "low";

dffeas \tdl_arr[2] (
	.clk(clk),
	.d(\tdl_arr[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[2]~q ),
	.prn(vcc));
defparam \tdl_arr[2] .is_wysiwyg = "true";
defparam \tdl_arr[2] .power_up = "low";

dffeas \tdl_arr[3] (
	.clk(clk),
	.d(\tdl_arr[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[3]~q ),
	.prn(vcc));
defparam \tdl_arr[3] .is_wysiwyg = "true";
defparam \tdl_arr[3] .power_up = "low";

dffeas \tdl_arr[4] (
	.clk(clk),
	.d(\tdl_arr[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\tdl_arr[4]~q ),
	.prn(vcc));
defparam \tdl_arr[4] .is_wysiwyg = "true";
defparam \tdl_arr[4] .power_up = "low";

endmodule

module IFFT_asj_fft_twadgen (
	global_clock_enable,
	twad_tdl_0_6,
	twad_tdl_1_6,
	twad_tdl_2_6,
	twad_tdl_3_6,
	Mux1,
	Mux0,
	Mux11,
	Mux01,
	clk)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	twad_tdl_0_6;
output 	twad_tdl_1_6;
output 	twad_tdl_2_6;
output 	twad_tdl_3_6;
input 	Mux1;
input 	Mux0;
input 	Mux11;
input 	Mux01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \twad_temp[0]~q ;
wire \twad_tdl[0][0]~q ;
wire \twad_tdl[1][0]~q ;
wire \twad_tdl[2][0]~q ;
wire \twad_tdl[3][0]~q ;
wire \twad_tdl[4][0]~q ;
wire \twad_tdl[5][0]~q ;
wire \twad_temp[1]~q ;
wire \twad_tdl[0][1]~q ;
wire \twad_tdl[1][1]~q ;
wire \twad_tdl[2][1]~q ;
wire \twad_tdl[3][1]~q ;
wire \twad_tdl[4][1]~q ;
wire \twad_tdl[5][1]~q ;
wire \twad_temp[2]~q ;
wire \twad_tdl[0][2]~q ;
wire \twad_tdl[1][2]~q ;
wire \twad_tdl[2][2]~q ;
wire \twad_tdl[3][2]~q ;
wire \twad_tdl[4][2]~q ;
wire \twad_tdl[5][2]~q ;
wire \twad_temp[3]~q ;
wire \twad_tdl[0][3]~q ;
wire \twad_tdl[1][3]~q ;
wire \twad_tdl[2][3]~q ;
wire \twad_tdl[3][3]~q ;
wire \twad_tdl[4][3]~q ;
wire \twad_tdl[5][3]~q ;


dffeas \twad_tdl[6][0] (
	.clk(clk),
	.d(\twad_tdl[5][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(twad_tdl_0_6),
	.prn(vcc));
defparam \twad_tdl[6][0] .is_wysiwyg = "true";
defparam \twad_tdl[6][0] .power_up = "low";

dffeas \twad_tdl[6][1] (
	.clk(clk),
	.d(\twad_tdl[5][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(twad_tdl_1_6),
	.prn(vcc));
defparam \twad_tdl[6][1] .is_wysiwyg = "true";
defparam \twad_tdl[6][1] .power_up = "low";

dffeas \twad_tdl[6][2] (
	.clk(clk),
	.d(\twad_tdl[5][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(twad_tdl_2_6),
	.prn(vcc));
defparam \twad_tdl[6][2] .is_wysiwyg = "true";
defparam \twad_tdl[6][2] .power_up = "low";

dffeas \twad_tdl[6][3] (
	.clk(clk),
	.d(\twad_tdl[5][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(twad_tdl_3_6),
	.prn(vcc));
defparam \twad_tdl[6][3] .is_wysiwyg = "true";
defparam \twad_tdl[6][3] .power_up = "low";

dffeas \twad_temp[0] (
	.clk(clk),
	.d(Mux1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_temp[0]~q ),
	.prn(vcc));
defparam \twad_temp[0] .is_wysiwyg = "true";
defparam \twad_temp[0] .power_up = "low";

dffeas \twad_tdl[0][0] (
	.clk(clk),
	.d(\twad_temp[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[0][0]~q ),
	.prn(vcc));
defparam \twad_tdl[0][0] .is_wysiwyg = "true";
defparam \twad_tdl[0][0] .power_up = "low";

dffeas \twad_tdl[1][0] (
	.clk(clk),
	.d(\twad_tdl[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[1][0]~q ),
	.prn(vcc));
defparam \twad_tdl[1][0] .is_wysiwyg = "true";
defparam \twad_tdl[1][0] .power_up = "low";

dffeas \twad_tdl[2][0] (
	.clk(clk),
	.d(\twad_tdl[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[2][0]~q ),
	.prn(vcc));
defparam \twad_tdl[2][0] .is_wysiwyg = "true";
defparam \twad_tdl[2][0] .power_up = "low";

dffeas \twad_tdl[3][0] (
	.clk(clk),
	.d(\twad_tdl[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[3][0]~q ),
	.prn(vcc));
defparam \twad_tdl[3][0] .is_wysiwyg = "true";
defparam \twad_tdl[3][0] .power_up = "low";

dffeas \twad_tdl[4][0] (
	.clk(clk),
	.d(\twad_tdl[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[4][0]~q ),
	.prn(vcc));
defparam \twad_tdl[4][0] .is_wysiwyg = "true";
defparam \twad_tdl[4][0] .power_up = "low";

dffeas \twad_tdl[5][0] (
	.clk(clk),
	.d(\twad_tdl[4][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[5][0]~q ),
	.prn(vcc));
defparam \twad_tdl[5][0] .is_wysiwyg = "true";
defparam \twad_tdl[5][0] .power_up = "low";

dffeas \twad_temp[1] (
	.clk(clk),
	.d(Mux0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_temp[1]~q ),
	.prn(vcc));
defparam \twad_temp[1] .is_wysiwyg = "true";
defparam \twad_temp[1] .power_up = "low";

dffeas \twad_tdl[0][1] (
	.clk(clk),
	.d(\twad_temp[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[0][1]~q ),
	.prn(vcc));
defparam \twad_tdl[0][1] .is_wysiwyg = "true";
defparam \twad_tdl[0][1] .power_up = "low";

dffeas \twad_tdl[1][1] (
	.clk(clk),
	.d(\twad_tdl[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[1][1]~q ),
	.prn(vcc));
defparam \twad_tdl[1][1] .is_wysiwyg = "true";
defparam \twad_tdl[1][1] .power_up = "low";

dffeas \twad_tdl[2][1] (
	.clk(clk),
	.d(\twad_tdl[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[2][1]~q ),
	.prn(vcc));
defparam \twad_tdl[2][1] .is_wysiwyg = "true";
defparam \twad_tdl[2][1] .power_up = "low";

dffeas \twad_tdl[3][1] (
	.clk(clk),
	.d(\twad_tdl[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[3][1]~q ),
	.prn(vcc));
defparam \twad_tdl[3][1] .is_wysiwyg = "true";
defparam \twad_tdl[3][1] .power_up = "low";

dffeas \twad_tdl[4][1] (
	.clk(clk),
	.d(\twad_tdl[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[4][1]~q ),
	.prn(vcc));
defparam \twad_tdl[4][1] .is_wysiwyg = "true";
defparam \twad_tdl[4][1] .power_up = "low";

dffeas \twad_tdl[5][1] (
	.clk(clk),
	.d(\twad_tdl[4][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[5][1]~q ),
	.prn(vcc));
defparam \twad_tdl[5][1] .is_wysiwyg = "true";
defparam \twad_tdl[5][1] .power_up = "low";

dffeas \twad_temp[2] (
	.clk(clk),
	.d(Mux11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_temp[2]~q ),
	.prn(vcc));
defparam \twad_temp[2] .is_wysiwyg = "true";
defparam \twad_temp[2] .power_up = "low";

dffeas \twad_tdl[0][2] (
	.clk(clk),
	.d(\twad_temp[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[0][2]~q ),
	.prn(vcc));
defparam \twad_tdl[0][2] .is_wysiwyg = "true";
defparam \twad_tdl[0][2] .power_up = "low";

dffeas \twad_tdl[1][2] (
	.clk(clk),
	.d(\twad_tdl[0][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[1][2]~q ),
	.prn(vcc));
defparam \twad_tdl[1][2] .is_wysiwyg = "true";
defparam \twad_tdl[1][2] .power_up = "low";

dffeas \twad_tdl[2][2] (
	.clk(clk),
	.d(\twad_tdl[1][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[2][2]~q ),
	.prn(vcc));
defparam \twad_tdl[2][2] .is_wysiwyg = "true";
defparam \twad_tdl[2][2] .power_up = "low";

dffeas \twad_tdl[3][2] (
	.clk(clk),
	.d(\twad_tdl[2][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[3][2]~q ),
	.prn(vcc));
defparam \twad_tdl[3][2] .is_wysiwyg = "true";
defparam \twad_tdl[3][2] .power_up = "low";

dffeas \twad_tdl[4][2] (
	.clk(clk),
	.d(\twad_tdl[3][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[4][2]~q ),
	.prn(vcc));
defparam \twad_tdl[4][2] .is_wysiwyg = "true";
defparam \twad_tdl[4][2] .power_up = "low";

dffeas \twad_tdl[5][2] (
	.clk(clk),
	.d(\twad_tdl[4][2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[5][2]~q ),
	.prn(vcc));
defparam \twad_tdl[5][2] .is_wysiwyg = "true";
defparam \twad_tdl[5][2] .power_up = "low";

dffeas \twad_temp[3] (
	.clk(clk),
	.d(Mux01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_temp[3]~q ),
	.prn(vcc));
defparam \twad_temp[3] .is_wysiwyg = "true";
defparam \twad_temp[3] .power_up = "low";

dffeas \twad_tdl[0][3] (
	.clk(clk),
	.d(\twad_temp[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[0][3]~q ),
	.prn(vcc));
defparam \twad_tdl[0][3] .is_wysiwyg = "true";
defparam \twad_tdl[0][3] .power_up = "low";

dffeas \twad_tdl[1][3] (
	.clk(clk),
	.d(\twad_tdl[0][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[1][3]~q ),
	.prn(vcc));
defparam \twad_tdl[1][3] .is_wysiwyg = "true";
defparam \twad_tdl[1][3] .power_up = "low";

dffeas \twad_tdl[2][3] (
	.clk(clk),
	.d(\twad_tdl[1][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[2][3]~q ),
	.prn(vcc));
defparam \twad_tdl[2][3] .is_wysiwyg = "true";
defparam \twad_tdl[2][3] .power_up = "low";

dffeas \twad_tdl[3][3] (
	.clk(clk),
	.d(\twad_tdl[2][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[3][3]~q ),
	.prn(vcc));
defparam \twad_tdl[3][3] .is_wysiwyg = "true";
defparam \twad_tdl[3][3] .power_up = "low";

dffeas \twad_tdl[4][3] (
	.clk(clk),
	.d(\twad_tdl[3][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[4][3]~q ),
	.prn(vcc));
defparam \twad_tdl[4][3] .is_wysiwyg = "true";
defparam \twad_tdl[4][3] .power_up = "low";

dffeas \twad_tdl[5][3] (
	.clk(clk),
	.d(\twad_tdl[4][3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\twad_tdl[5][3]~q ),
	.prn(vcc));
defparam \twad_tdl[5][3] .is_wysiwyg = "true";
defparam \twad_tdl[5][3] .power_up = "low";

endmodule

module IFFT_asj_fft_wrengen (
	global_clock_enable,
	wc_i1,
	wd_i1,
	ram_a_not_b_vec_26,
	p_cd_en_0,
	p_cd_en_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	global_clock_enable;
output 	wc_i1;
output 	wd_i1;
input 	ram_a_not_b_vec_26;
input 	p_cd_en_0;
input 	p_cd_en_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wc_i~0_combout ;
wire \wd_i~0_combout ;


dffeas wc_i(
	.clk(clk),
	.d(\wc_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wc_i1),
	.prn(vcc));
defparam wc_i.is_wysiwyg = "true";
defparam wc_i.power_up = "low";

dffeas wd_i(
	.clk(clk),
	.d(\wd_i~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(wd_i1),
	.prn(vcc));
defparam wd_i.is_wysiwyg = "true";
defparam wd_i.power_up = "low";

cyclonev_lcell_comb \wc_i~0 (
	.dataa(!reset_n),
	.datab(!ram_a_not_b_vec_26),
	.datac(!p_cd_en_0),
	.datad(!p_cd_en_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wc_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wc_i~0 .extended_lut = "off";
defparam \wc_i~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \wc_i~0 .shared_arith = "off";

cyclonev_lcell_comb \wd_i~0 (
	.dataa(!reset_n),
	.datab(!ram_a_not_b_vec_26),
	.datac(!p_cd_en_0),
	.datad(!p_cd_en_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wd_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wd_i~0 .extended_lut = "off";
defparam \wd_i~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \wd_i~0 .shared_arith = "off";

endmodule

module IFFT_asj_fft_wrswgen (
	ram_block6a3,
	ram_block6a2,
	ram_block6a0,
	ram_block6a1,
	global_clock_enable,
	p_tdl_0_0,
	p_tdl_1_0,
	k_count_1,
	k_count_3,
	k_count_0,
	k_count_2,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ram_block6a3;
output 	ram_block6a2;
output 	ram_block6a0;
output 	ram_block6a1;
input 	global_clock_enable;
input 	p_tdl_0_0;
input 	p_tdl_1_0;
input 	k_count_1;
input 	k_count_3;
input 	k_count_0;
input 	k_count_2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux0~0_combout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ;
wire \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ;
wire \swa_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \swa_rtl_0|auto_generated|op_1~1_sumout ;
wire \swa_rtl_0|auto_generated|dffe3a[0]~q ;
wire \swa_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ;
wire \swa_rtl_0|auto_generated|op_1~2 ;
wire \swa_rtl_0|auto_generated|op_1~5_sumout ;
wire \swa_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \swa_rtl_0|auto_generated|dffe3a[1]~q ;
wire \swa_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \swa_rtl_0|auto_generated|op_1~6 ;
wire \swa_rtl_0|auto_generated|op_1~9_sumout ;
wire \swa_rtl_0|auto_generated|dffe3a[2]~q ;
wire \swa_rtl_0|auto_generated|op_1~10 ;
wire \swa_rtl_0|auto_generated|op_1~13_sumout ;
wire \swa_rtl_0|auto_generated|dffe3a[3]~q ;
wire \swa_rtl_0|auto_generated|op_1~14 ;
wire \swa_rtl_0|auto_generated|op_1~17_sumout ;
wire \swa_rtl_0|auto_generated|dffe3a[4]~q ;
wire \Mux1~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;

wire [143:0] \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3_PORTBDATAOUT_bus ;
wire [143:0] \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2_PORTBDATAOUT_bus ;
wire [143:0] \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0_PORTBDATAOUT_bus ;
wire [143:0] \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1_PORTBDATAOUT_bus ;

assign ram_block6a3 = \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3_PORTBDATAOUT_bus [0];

assign ram_block6a2 = \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2_PORTBDATAOUT_bus [0];

assign ram_block6a0 = \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0_PORTBDATAOUT_bus [0];

assign ram_block6a1 = \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1_PORTBDATAOUT_bus [0];

cyclonev_ram_block \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux0~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|dffe3a[4]~q ,\swa_rtl_0|auto_generated|dffe3a[3]~q ,\swa_rtl_0|auto_generated|dffe3a[2]~q ,\swa_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\swa_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\swa_rtl_0|auto_generated|altsyncram5|ram_block6a3_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .clk0_core_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .clk0_input_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .clk1_output_clock_enable = "ena1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .data_interleave_offset_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .data_interleave_width_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_wrswgen:\\gen_wrsw_1:get_wr_swtiches|altshift_taps:swa_rtl_0|shift_taps_dgv:auto_generated|altsyncram_vr91:altsyncram5|ALTSYNCRAM";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .mixed_port_feed_through_mode = "dont_care";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .operation_mode = "dual_port";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_data_out_clock = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_first_bit_number = 3;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_address_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_data_out_clock = "clock1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_first_bit_number = 3;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .port_b_read_enable_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a3 .ram_block_type = "auto";

cyclonev_ram_block \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux1~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|dffe3a[4]~q ,\swa_rtl_0|auto_generated|dffe3a[3]~q ,\swa_rtl_0|auto_generated|dffe3a[2]~q ,\swa_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\swa_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\swa_rtl_0|auto_generated|altsyncram5|ram_block6a2_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .clk0_core_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .clk0_input_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .clk1_output_clock_enable = "ena1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .data_interleave_offset_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .data_interleave_width_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_wrswgen:\\gen_wrsw_1:get_wr_swtiches|altshift_taps:swa_rtl_0|shift_taps_dgv:auto_generated|altsyncram_vr91:altsyncram5|ALTSYNCRAM";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .mixed_port_feed_through_mode = "dont_care";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .operation_mode = "dual_port";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_data_out_clock = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_first_bit_number = 2;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_address_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_data_out_clock = "clock1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_first_bit_number = 2;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .port_b_read_enable_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a2 .ram_block_type = "auto";

cyclonev_ram_block \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux3~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|dffe3a[4]~q ,\swa_rtl_0|auto_generated|dffe3a[3]~q ,\swa_rtl_0|auto_generated|dffe3a[2]~q ,\swa_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\swa_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\swa_rtl_0|auto_generated|altsyncram5|ram_block6a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .clk0_core_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .clk0_input_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .clk1_output_clock_enable = "ena1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .data_interleave_offset_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .data_interleave_width_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_wrswgen:\\gen_wrsw_1:get_wr_swtiches|altshift_taps:swa_rtl_0|shift_taps_dgv:auto_generated|altsyncram_vr91:altsyncram5|ALTSYNCRAM";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .mixed_port_feed_through_mode = "dont_care";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .operation_mode = "dual_port";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_data_out_clock = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_first_bit_number = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_address_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_data_out_clock = "clock1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_first_bit_number = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .port_b_read_enable_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a0 .ram_block_type = "auto";

cyclonev_ram_block \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(!global_clock_enable),
	.ena1(!global_clock_enable),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\Mux2~0_combout }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\swa_rtl_0|auto_generated|dffe3a[4]~q ,\swa_rtl_0|auto_generated|dffe3a[3]~q ,\swa_rtl_0|auto_generated|dffe3a[2]~q ,\swa_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\swa_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\swa_rtl_0|auto_generated|altsyncram5|ram_block6a1_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .clk0_core_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .clk0_input_clock_enable = "ena0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .clk1_output_clock_enable = "ena1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .data_interleave_offset_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .data_interleave_width_in_bits = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|asj_fft_wrswgen:\\gen_wrsw_1:get_wr_swtiches|altshift_taps:swa_rtl_0|shift_taps_dgv:auto_generated|altsyncram_vr91:altsyncram5|ALTSYNCRAM";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .mixed_port_feed_through_mode = "dont_care";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .operation_mode = "dual_port";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_data_out_clock = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_first_bit_number = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_address_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_address_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_address_width = 5;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_data_out_clear = "none";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_data_out_clock = "clock1";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_data_width = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_first_address = 0;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_first_bit_number = 1;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_last_address = 17;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_logical_ram_depth = 18;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_logical_ram_width = 4;
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .port_b_read_enable_clock = "clock0";
defparam \swa_rtl_0|auto_generated|altsyncram5|ram_block6a1 .ram_block_type = "auto";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!p_tdl_0_0),
	.datab(!p_tdl_1_0),
	.datac(!k_count_1),
	.datad(!k_count_3),
	.datae(!k_count_0),
	.dataf(!k_count_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h6996966996696996;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\swa_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\swa_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\swa_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.cout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\swa_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ),
	.cout(),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .lut_mask = 64'h0000000000000000;
defparam \swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .shared_arith = "off";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(!\swa_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\swa_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \swa_rtl_0|auto_generated|cntr1|cout_actual .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \swa_rtl_0|auto_generated|cntr1|cout_actual .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\swa_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\swa_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \swa_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|dffe3a[0] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|cmpr4_aeb_int~0 (
	.dataa(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\swa_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \swa_rtl_0|auto_generated|cmpr4_aeb_int~0 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|cmpr4_aeb_int~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \swa_rtl_0|auto_generated|cmpr4_aeb_int~0 .shared_arith = "off";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|op_1~5 (
	.dataa(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(!\swa_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\swa_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \swa_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h000055FF000000FF;
defparam \swa_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\swa_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\swa_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \swa_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \swa_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|dffe3a[1] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\swa_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\swa_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \swa_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \swa_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\swa_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \swa_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|dffe3a[2] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(\swa_rtl_0|auto_generated|op_1~14 ),
	.shareout());
defparam \swa_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \swa_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|dffe3a[3] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_lcell_comb \swa_rtl_0|auto_generated|op_1~17 (
	.dataa(!\swa_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\swa_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\swa_rtl_0|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\swa_rtl_0|auto_generated|op_1~17_sumout ),
	.cout(),
	.shareout());
defparam \swa_rtl_0|auto_generated|op_1~17 .extended_lut = "off";
defparam \swa_rtl_0|auto_generated|op_1~17 .lut_mask = 64'h0000FFAA00005555;
defparam \swa_rtl_0|auto_generated|op_1~17 .shared_arith = "off";

dffeas \swa_rtl_0|auto_generated|dffe3a[4] (
	.clk(clk),
	.d(\swa_rtl_0|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!global_clock_enable),
	.q(\swa_rtl_0|auto_generated|dffe3a[4]~q ),
	.prn(vcc));
defparam \swa_rtl_0|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \swa_rtl_0|auto_generated|dffe3a[4] .power_up = "low";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!p_tdl_0_0),
	.datab(!p_tdl_1_0),
	.datac(!k_count_0),
	.datad(!k_count_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h6996699669966996;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!p_tdl_0_0),
	.datab(!p_tdl_1_0),
	.datac(!k_count_0),
	.datad(!k_count_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!p_tdl_0_0),
	.datab(!p_tdl_1_0),
	.datac(!k_count_1),
	.datad(!k_count_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \Mux2~0 .shared_arith = "off";

endmodule

module IFFT_auk_dspip_avalon_streaming_controller (
	sink_in_work,
	at_source_valid_s,
	source_packet_error_1,
	source_packet_error_0,
	sink_stall,
	sink_stall_reg1,
	source_stall_reg1,
	sink_ready_ctrl,
	master_sink_ena,
	send_eop_s,
	packet_error_s_1,
	packet_error_s_0,
	stall_controller_comb,
	stall_reg1,
	sink_ready_ctrl1,
	Mux0,
	Mux01,
	Mux02,
	stall_controller_comb1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sink_in_work;
input 	at_source_valid_s;
output 	source_packet_error_1;
output 	source_packet_error_0;
input 	sink_stall;
output 	sink_stall_reg1;
output 	source_stall_reg1;
output 	sink_ready_ctrl;
input 	master_sink_ena;
input 	send_eop_s;
input 	packet_error_s_1;
input 	packet_error_s_0;
input 	stall_controller_comb;
output 	stall_reg1;
output 	sink_ready_ctrl1;
input 	Mux0;
input 	Mux01;
input 	Mux02;
input 	stall_controller_comb1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_stall_reg~0_combout ;
wire \source_stall_reg~0_combout ;
wire \stall_int~combout ;


dffeas \source_packet_error[1] (
	.clk(clk),
	.d(packet_error_s_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_1),
	.prn(vcc));
defparam \source_packet_error[1] .is_wysiwyg = "true";
defparam \source_packet_error[1] .power_up = "low";

dffeas \source_packet_error[0] (
	.clk(clk),
	.d(packet_error_s_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_packet_error_0),
	.prn(vcc));
defparam \source_packet_error[0] .is_wysiwyg = "true";
defparam \source_packet_error[0] .power_up = "low";

dffeas sink_stall_reg(
	.clk(clk),
	.d(\sink_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sink_stall_reg1),
	.prn(vcc));
defparam sink_stall_reg.is_wysiwyg = "true";
defparam sink_stall_reg.power_up = "low";

dffeas source_stall_reg(
	.clk(clk),
	.d(\source_stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_reg1),
	.prn(vcc));
defparam source_stall_reg.is_wysiwyg = "true";
defparam source_stall_reg.power_up = "low";

cyclonev_lcell_comb \sink_ready_ctrl~0 (
	.dataa(!sink_stall_reg1),
	.datab(!source_stall_reg1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready_ctrl),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready_ctrl~0 .extended_lut = "off";
defparam \sink_ready_ctrl~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \sink_ready_ctrl~0 .shared_arith = "off";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_int~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

cyclonev_lcell_comb \sink_ready_ctrl~1 (
	.dataa(!sink_stall_reg1),
	.datab(!source_stall_reg1),
	.datac(!master_sink_ena),
	.datad(!send_eop_s),
	.datae(!sink_in_work),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready_ctrl1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready_ctrl~1 .extended_lut = "off";
defparam \sink_ready_ctrl~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \sink_ready_ctrl~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_stall_reg~0 (
	.dataa(!sink_stall),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_stall_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_stall_reg~0 .extended_lut = "off";
defparam \sink_stall_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sink_stall_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \source_stall_reg~0 (
	.dataa(!Mux02),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_stall_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_stall_reg~0 .extended_lut = "off";
defparam \source_stall_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \source_stall_reg~0 .shared_arith = "off";

cyclonev_lcell_comb stall_int(
	.dataa(!at_source_valid_s),
	.datab(!sink_stall),
	.datac(!stall_controller_comb),
	.datad(!stall_controller_comb1),
	.datae(!Mux0),
	.dataf(!Mux01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stall_int~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam stall_int.extended_lut = "off";
defparam stall_int.lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam stall_int.shared_arith = "off";

endmodule

module IFFT_auk_dspip_avalon_streaming_sink (
	sink_in_work,
	q_b_14,
	q_b_6,
	q_b_13,
	q_b_5,
	q_b_10,
	q_b_2,
	q_b_11,
	q_b_3,
	q_b_12,
	q_b_4,
	q_b_15,
	q_b_7,
	q_b_8,
	q_b_0,
	q_b_9,
	q_b_1,
	at_sink_ready_s1,
	sink_stall1,
	sink_stall_reg,
	source_stall_reg,
	sink_ready_ctrl,
	master_sink_ena,
	send_eop_s1,
	packet_error_s_1,
	packet_error_s_0,
	send_sop_s1,
	sink_ready_ctrl1,
	clk,
	reset_n,
	sink_eop,
	sink_valid,
	sink_error_0,
	sink_error_1,
	sink_sop,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
input 	sink_in_work;
output 	q_b_14;
output 	q_b_6;
output 	q_b_13;
output 	q_b_5;
output 	q_b_10;
output 	q_b_2;
output 	q_b_11;
output 	q_b_3;
output 	q_b_12;
output 	q_b_4;
output 	q_b_15;
output 	q_b_7;
output 	q_b_8;
output 	q_b_0;
output 	q_b_9;
output 	q_b_1;
output 	at_sink_ready_s1;
output 	sink_stall1;
input 	sink_stall_reg;
input 	source_stall_reg;
input 	sink_ready_ctrl;
input 	master_sink_ena;
output 	send_eop_s1;
output 	packet_error_s_1;
output 	packet_error_s_0;
output 	send_sop_s1;
input 	sink_ready_ctrl1;
input 	clk;
input 	reset_n;
input 	sink_eop;
input 	sink_valid;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_sop;
input 	[15:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \fifo_wrreq~0_combout ;
wire \at_sink_data_int[14]~q ;
wire \at_sink_data_int[6]~q ;
wire \at_sink_data_int[13]~q ;
wire \at_sink_data_int[5]~q ;
wire \at_sink_data_int[10]~q ;
wire \at_sink_data_int[2]~q ;
wire \at_sink_data_int[11]~q ;
wire \at_sink_data_int[3]~q ;
wire \at_sink_data_int[12]~q ;
wire \at_sink_data_int[4]~q ;
wire \at_sink_data_int[15]~q ;
wire \at_sink_data_int[7]~q ;
wire \at_sink_data_int[8]~q ;
wire \at_sink_data_int[0]~q ;
wire \at_sink_data_int[9]~q ;
wire \at_sink_data_int[1]~q ;
wire \data_take~combout ;
wire \at_sink_ready_s~0_combout ;
wire \sink_start~0_combout ;
wire \sink_start~q ;
wire \out_cnt[0]~6_combout ;
wire \Selector7~2_combout ;
wire \sink_stall_s~q ;
wire \Selector8~0_combout ;
wire \sink_out_state.normal~q ;
wire \Selector10~0_combout ;
wire \sink_out_state.empty_and_ready~q ;
wire \Selector7~3_combout ;
wire \out_cnt[0]~q ;
wire \out_cnt~4_combout ;
wire \out_cnt[1]~q ;
wire \out_cnt~3_combout ;
wire \out_cnt[2]~q ;
wire \out_cnt~2_combout ;
wire \out_cnt[3]~q ;
wire \Equal2~0_combout ;
wire \out_cnt~1_combout ;
wire \out_cnt[4]~q ;
wire \out_cnt~0_combout ;
wire \out_cnt[5]~q ;
wire \Equal2~1_combout ;
wire \send_sop_eop_p~0_combout ;
wire \at_sink_error_int~0_combout ;
wire \sink_comb_update_2~0_combout ;
wire \Selector3~6_combout ;
wire \Selector3~7_combout ;
wire \Selector3~3_combout ;
wire \Selector3~8_combout ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \Selector3~2_combout ;
wire \Selector3~5_combout ;
wire \sink_state.st_err~q ;
wire \Selector3~4_combout ;
wire \count~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~6_combout ;
wire \Selector2~4_combout ;
wire \Selector2~2_combout ;
wire \Selector4~1_combout ;
wire \Selector4~0_combout ;
wire \count[0]~1_combout ;
wire \count[0]~q ;
wire \count~5_combout ;
wire \count[1]~q ;
wire \count~6_combout ;
wire \count[2]~q ;
wire \Add0~2_combout ;
wire \count~4_combout ;
wire \count[3]~q ;
wire \Add0~1_combout ;
wire \count~3_combout ;
wire \count[4]~q ;
wire \Add0~0_combout ;
wire \count~2_combout ;
wire \count[5]~q ;
wire \max_reached~0_combout ;
wire \max_reached~1_combout ;
wire \max_reached~q ;
wire \Selector2~5_combout ;
wire \Selector2~3_combout ;
wire \sink_state.run1~q ;
wire \Selector2~0_combout ;
wire \Selector1~0_combout ;
wire \sink_state.stall~q ;
wire \packet_error_int~0_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \sink_state.end1~q ;
wire \Selector0~0_combout ;
wire \sink_state.start~q ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \Equal1~0_combout ;


IFFT_scfifo_1 \normal_fifo:fifo_eab_on:in_fifo (
	.q({q_unconnected_wire_17,q_unconnected_wire_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.dffe_af(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.counter_reg_bit_0(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.empty_dff(\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.sink_out_stateempty_and_ready(\sink_out_state.empty_and_ready~q ),
	.Selector7(\Selector7~0_combout ),
	.sink_stall(sink_stall1),
	.Selector71(\Selector7~1_combout ),
	.wrreq(\fifo_wrreq~0_combout ),
	.Selector72(\Selector7~2_combout ),
	.out_cnt_0(\out_cnt[0]~q ),
	.rdreq(\Selector7~3_combout ),
	.data({gnd,gnd,\at_sink_data_int[15]~q ,\at_sink_data_int[14]~q ,\at_sink_data_int[13]~q ,\at_sink_data_int[12]~q ,\at_sink_data_int[11]~q ,\at_sink_data_int[10]~q ,\at_sink_data_int[9]~q ,\at_sink_data_int[8]~q ,\at_sink_data_int[7]~q ,\at_sink_data_int[6]~q ,
\at_sink_data_int[5]~q ,\at_sink_data_int[4]~q ,\at_sink_data_int[3]~q ,\at_sink_data_int[2]~q ,\at_sink_data_int[1]~q ,\at_sink_data_int[0]~q }),
	.clock(clk),
	.reset_n(reset_n));

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!\sink_start~q ),
	.datab(!\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.datac(!\sink_out_state.empty_and_ready~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector7~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~1 (
	.dataa(!sink_stall1),
	.datab(!\sink_out_state.normal~q ),
	.datac(!sink_ready_ctrl),
	.datad(!master_sink_ena),
	.datae(!send_eop_s1),
	.dataf(!sink_in_work),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~1 .extended_lut = "off";
defparam \Selector7~1 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Selector7~1 .shared_arith = "off";

cyclonev_lcell_comb \fifo_wrreq~0 (
	.dataa(!\sink_state.run1~q ),
	.datab(!\sink_state.end1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wrreq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wrreq~0 .extended_lut = "off";
defparam \fifo_wrreq~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \fifo_wrreq~0 .shared_arith = "off";

dffeas \at_sink_data_int[14] (
	.clk(clk),
	.d(at_sink_data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[14]~q ),
	.prn(vcc));
defparam \at_sink_data_int[14] .is_wysiwyg = "true";
defparam \at_sink_data_int[14] .power_up = "low";

dffeas \at_sink_data_int[6] (
	.clk(clk),
	.d(at_sink_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[6]~q ),
	.prn(vcc));
defparam \at_sink_data_int[6] .is_wysiwyg = "true";
defparam \at_sink_data_int[6] .power_up = "low";

dffeas \at_sink_data_int[13] (
	.clk(clk),
	.d(at_sink_data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[13]~q ),
	.prn(vcc));
defparam \at_sink_data_int[13] .is_wysiwyg = "true";
defparam \at_sink_data_int[13] .power_up = "low";

dffeas \at_sink_data_int[5] (
	.clk(clk),
	.d(at_sink_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[5]~q ),
	.prn(vcc));
defparam \at_sink_data_int[5] .is_wysiwyg = "true";
defparam \at_sink_data_int[5] .power_up = "low";

dffeas \at_sink_data_int[10] (
	.clk(clk),
	.d(at_sink_data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[10]~q ),
	.prn(vcc));
defparam \at_sink_data_int[10] .is_wysiwyg = "true";
defparam \at_sink_data_int[10] .power_up = "low";

dffeas \at_sink_data_int[2] (
	.clk(clk),
	.d(at_sink_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[2]~q ),
	.prn(vcc));
defparam \at_sink_data_int[2] .is_wysiwyg = "true";
defparam \at_sink_data_int[2] .power_up = "low";

dffeas \at_sink_data_int[11] (
	.clk(clk),
	.d(at_sink_data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[11]~q ),
	.prn(vcc));
defparam \at_sink_data_int[11] .is_wysiwyg = "true";
defparam \at_sink_data_int[11] .power_up = "low";

dffeas \at_sink_data_int[3] (
	.clk(clk),
	.d(at_sink_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[3]~q ),
	.prn(vcc));
defparam \at_sink_data_int[3] .is_wysiwyg = "true";
defparam \at_sink_data_int[3] .power_up = "low";

dffeas \at_sink_data_int[12] (
	.clk(clk),
	.d(at_sink_data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[12]~q ),
	.prn(vcc));
defparam \at_sink_data_int[12] .is_wysiwyg = "true";
defparam \at_sink_data_int[12] .power_up = "low";

dffeas \at_sink_data_int[4] (
	.clk(clk),
	.d(at_sink_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[4]~q ),
	.prn(vcc));
defparam \at_sink_data_int[4] .is_wysiwyg = "true";
defparam \at_sink_data_int[4] .power_up = "low";

dffeas \at_sink_data_int[15] (
	.clk(clk),
	.d(at_sink_data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[15]~q ),
	.prn(vcc));
defparam \at_sink_data_int[15] .is_wysiwyg = "true";
defparam \at_sink_data_int[15] .power_up = "low";

dffeas \at_sink_data_int[7] (
	.clk(clk),
	.d(at_sink_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[7]~q ),
	.prn(vcc));
defparam \at_sink_data_int[7] .is_wysiwyg = "true";
defparam \at_sink_data_int[7] .power_up = "low";

dffeas \at_sink_data_int[8] (
	.clk(clk),
	.d(at_sink_data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[8]~q ),
	.prn(vcc));
defparam \at_sink_data_int[8] .is_wysiwyg = "true";
defparam \at_sink_data_int[8] .power_up = "low";

dffeas \at_sink_data_int[0] (
	.clk(clk),
	.d(at_sink_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[0]~q ),
	.prn(vcc));
defparam \at_sink_data_int[0] .is_wysiwyg = "true";
defparam \at_sink_data_int[0] .power_up = "low";

dffeas \at_sink_data_int[9] (
	.clk(clk),
	.d(at_sink_data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[9]~q ),
	.prn(vcc));
defparam \at_sink_data_int[9] .is_wysiwyg = "true";
defparam \at_sink_data_int[9] .power_up = "low";

dffeas \at_sink_data_int[1] (
	.clk(clk),
	.d(at_sink_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data_take~combout ),
	.q(\at_sink_data_int[1]~q ),
	.prn(vcc));
defparam \at_sink_data_int[1] .is_wysiwyg = "true";
defparam \at_sink_data_int[1] .power_up = "low";

cyclonev_lcell_comb data_take(
	.dataa(!\fifo_wrreq~0_combout ),
	.datab(!\Selector3~6_combout ),
	.datac(!\Selector2~4_combout ),
	.datad(!\Selector2~2_combout ),
	.datae(!\Selector4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_take~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam data_take.extended_lut = "off";
defparam data_take.lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam data_take.shared_arith = "off";

dffeas at_sink_ready_s(
	.clk(clk),
	.d(\at_sink_ready_s~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_sink_ready_s1),
	.prn(vcc));
defparam at_sink_ready_s.is_wysiwyg = "true";
defparam at_sink_ready_s.power_up = "low";

cyclonev_lcell_comb sink_stall(
	.dataa(!\sink_start~q ),
	.datab(!\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|empty_dff~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_stall1),
	.sumout(),
	.cout(),
	.shareout());
defparam sink_stall.extended_lut = "off";
defparam sink_stall.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam sink_stall.shared_arith = "off";

dffeas send_eop_s(
	.clk(clk),
	.d(\Equal2~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_eop_s1),
	.prn(vcc));
defparam send_eop_s.is_wysiwyg = "true";
defparam send_eop_s.power_up = "low";

dffeas \packet_error_s[1] (
	.clk(clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_1),
	.prn(vcc));
defparam \packet_error_s[1] .is_wysiwyg = "true";
defparam \packet_error_s[1] .power_up = "low";

dffeas \packet_error_s[0] (
	.clk(clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_error_s_0),
	.prn(vcc));
defparam \packet_error_s[0] .is_wysiwyg = "true";
defparam \packet_error_s[0] .power_up = "low";

dffeas send_sop_s(
	.clk(clk),
	.d(\Equal1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\send_sop_eop_p~0_combout ),
	.q(send_sop_s1),
	.prn(vcc));
defparam send_sop_s.is_wysiwyg = "true";
defparam send_sop_s.power_up = "low";

cyclonev_lcell_comb \at_sink_ready_s~0 (
	.dataa(!\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dffe_af~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\at_sink_ready_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \at_sink_ready_s~0 .extended_lut = "off";
defparam \at_sink_ready_s~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \at_sink_ready_s~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_start~0 (
	.dataa(!\normal_fifo:fifo_eab_on:in_fifo|auto_generated|dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(!\sink_start~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_start~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_start~0 .extended_lut = "off";
defparam \sink_start~0 .lut_mask = 64'h7777777777777777;
defparam \sink_start~0 .shared_arith = "off";

dffeas sink_start(
	.clk(clk),
	.d(\sink_start~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_start~q ),
	.prn(vcc));
defparam sink_start.is_wysiwyg = "true";
defparam sink_start.power_up = "low";

cyclonev_lcell_comb \out_cnt[0]~6 (
	.dataa(!\out_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cnt[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cnt[0]~6 .extended_lut = "off";
defparam \out_cnt[0]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \out_cnt[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~2 (
	.dataa(!\sink_out_state.normal~q ),
	.datab(!sink_stall_reg),
	.datac(!source_stall_reg),
	.datad(!master_sink_ena),
	.datae(!send_eop_s1),
	.dataf(!sink_in_work),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~2 .extended_lut = "off";
defparam \Selector7~2 .lut_mask = 64'hFFFFEFFFFFFFFFFF;
defparam \Selector7~2 .shared_arith = "off";

dffeas sink_stall_s(
	.clk(clk),
	.d(sink_stall1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_stall_s~q ),
	.prn(vcc));
defparam sink_stall_s.is_wysiwyg = "true";
defparam sink_stall_s.power_up = "low";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!sink_stall1),
	.datab(!\Selector7~2_combout ),
	.datac(!\sink_stall_s~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Selector8~0 .shared_arith = "off";

dffeas \sink_out_state.normal (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.normal~q ),
	.prn(vcc));
defparam \sink_out_state.normal .is_wysiwyg = "true";
defparam \sink_out_state.normal .power_up = "low";

cyclonev_lcell_comb \Selector10~0 (
	.dataa(!sink_stall1),
	.datab(!\sink_out_state.empty_and_ready~q ),
	.datac(!\sink_out_state.normal~q ),
	.datad(!sink_ready_ctrl1),
	.datae(!\sink_stall_s~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'hF7FFFFF7F7FFFFF7;
defparam \Selector10~0 .shared_arith = "off";

dffeas \sink_out_state.empty_and_ready (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_out_state.empty_and_ready~q ),
	.prn(vcc));
defparam \sink_out_state.empty_and_ready .is_wysiwyg = "true";
defparam \sink_out_state.empty_and_ready .power_up = "low";

cyclonev_lcell_comb \Selector7~3 (
	.dataa(!sink_stall1),
	.datab(!\sink_out_state.empty_and_ready~q ),
	.datac(!\Selector7~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~3 .extended_lut = "off";
defparam \Selector7~3 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Selector7~3 .shared_arith = "off";

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector7~3_combout ),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

cyclonev_lcell_comb \out_cnt~4 (
	.dataa(!\out_cnt[0]~q ),
	.datab(!\out_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cnt~4 .extended_lut = "off";
defparam \out_cnt~4 .lut_mask = 64'h6666666666666666;
defparam \out_cnt~4 .shared_arith = "off";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector7~3_combout ),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

cyclonev_lcell_comb \out_cnt~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\out_cnt[2]~q ),
	.datae(!\out_cnt[1]~q ),
	.dataf(!\out_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cnt~3 .extended_lut = "off";
defparam \out_cnt~3 .lut_mask = 64'hFF0000FF00FFFF00;
defparam \out_cnt~3 .shared_arith = "off";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector7~3_combout ),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

cyclonev_lcell_comb \out_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\out_cnt[3]~q ),
	.datad(!\out_cnt[2]~q ),
	.datae(!\out_cnt[1]~q ),
	.dataf(!\out_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cnt~2 .extended_lut = "off";
defparam \out_cnt~2 .lut_mask = 64'h0FF0F00FF00F0FF0;
defparam \out_cnt~2 .shared_arith = "off";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector7~3_combout ),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\out_cnt[3]~q ),
	.datab(!\out_cnt[2]~q ),
	.datac(!\out_cnt[1]~q ),
	.datad(!\out_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \out_cnt~1 (
	.dataa(gnd),
	.datab(!\out_cnt[4]~q ),
	.datac(!\Equal2~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cnt~1 .extended_lut = "off";
defparam \out_cnt~1 .lut_mask = 64'h3C3C3C3C3C3C3C3C;
defparam \out_cnt~1 .shared_arith = "off";

dffeas \out_cnt[4] (
	.clk(clk),
	.d(\out_cnt~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector7~3_combout ),
	.q(\out_cnt[4]~q ),
	.prn(vcc));
defparam \out_cnt[4] .is_wysiwyg = "true";
defparam \out_cnt[4] .power_up = "low";

cyclonev_lcell_comb \out_cnt~0 (
	.dataa(!\out_cnt[5]~q ),
	.datab(!\out_cnt[4]~q ),
	.datac(!\Equal2~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cnt~0 .extended_lut = "off";
defparam \out_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \out_cnt~0 .shared_arith = "off";

dffeas \out_cnt[5] (
	.clk(clk),
	.d(\out_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector7~3_combout ),
	.q(\out_cnt[5]~q ),
	.prn(vcc));
defparam \out_cnt[5] .is_wysiwyg = "true";
defparam \out_cnt[5] .power_up = "low";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!\out_cnt[5]~q ),
	.datab(!\out_cnt[4]~q ),
	.datac(!\Equal2~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \send_sop_eop_p~0 (
	.dataa(!sink_stall1),
	.datab(!\sink_out_state.empty_and_ready~q ),
	.datac(!\sink_out_state.normal~q ),
	.datad(!sink_ready_ctrl1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\send_sop_eop_p~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \send_sop_eop_p~0 .extended_lut = "off";
defparam \send_sop_eop_p~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \send_sop_eop_p~0 .shared_arith = "off";

cyclonev_lcell_comb \at_sink_error_int~0 (
	.dataa(!at_sink_ready_s1),
	.datab(!sink_valid),
	.datac(!sink_error_0),
	.datad(!sink_error_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\at_sink_error_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \at_sink_error_int~0 .extended_lut = "off";
defparam \at_sink_error_int~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \at_sink_error_int~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_comb_update_2~0 (
	.dataa(!at_sink_ready_s1),
	.datab(!sink_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_comb_update_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_comb_update_2~0 .extended_lut = "off";
defparam \sink_comb_update_2~0 .lut_mask = 64'h7777777777777777;
defparam \sink_comb_update_2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~6 (
	.dataa(!\sink_state.run1~q ),
	.datab(!\sink_state.stall~q ),
	.datac(!at_sink_ready_s1),
	.datad(!sink_valid),
	.datae(!sink_error_0),
	.dataf(!sink_error_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~6 .extended_lut = "off";
defparam \Selector3~6 .lut_mask = 64'h5F3FFFFFFFFFFFFF;
defparam \Selector3~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~7 (
	.dataa(!\max_reached~q ),
	.datab(!sink_eop),
	.datac(!sink_error_1),
	.datad(!sink_sop),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~7 .extended_lut = "off";
defparam \Selector3~7 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \Selector3~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~3 (
	.dataa(!\sink_state.run1~q ),
	.datab(!at_sink_ready_s1),
	.datac(!sink_valid),
	.datad(!sink_error_0),
	.datae(!\sink_state.stall~q ),
	.dataf(!\Selector3~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~3 .extended_lut = "off";
defparam \Selector3~3 .lut_mask = 64'hFFFFFFFFBFFF8FFF;
defparam \Selector3~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~8 (
	.dataa(!sink_error_0),
	.datab(!sink_error_1),
	.datac(!sink_sop),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~8 .extended_lut = "off";
defparam \Selector3~8 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Selector3~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!at_sink_ready_s1),
	.datab(!\max_reached~q ),
	.datac(!sink_eop),
	.datad(!sink_valid),
	.datae(!\sink_state.stall~q ),
	.dataf(!\Selector3~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!\sink_state.run1~q ),
	.datab(!\max_reached~q ),
	.datac(!sink_eop),
	.datad(!at_sink_ready_s1),
	.datae(!sink_valid),
	.dataf(!\Selector3~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \Selector3~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~2 (
	.dataa(!at_sink_ready_s1),
	.datab(!\max_reached~q ),
	.datac(!sink_eop),
	.datad(!sink_valid),
	.datae(!\at_sink_error_int~0_combout ),
	.dataf(!\Selector2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~2 .extended_lut = "off";
defparam \Selector3~2 .lut_mask = 64'hF3FFFFFF77FFFFFF;
defparam \Selector3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~5 (
	.dataa(!\Selector3~0_combout ),
	.datab(!\Selector3~1_combout ),
	.datac(!\Selector3~2_combout ),
	.datad(!\Selector3~3_combout ),
	.datae(!\Selector3~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~5 .extended_lut = "off";
defparam \Selector3~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector3~5 .shared_arith = "off";

dffeas \sink_state.st_err (
	.clk(clk),
	.d(\Selector3~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.st_err~q ),
	.prn(vcc));
defparam \sink_state.st_err .is_wysiwyg = "true";
defparam \sink_state.st_err .power_up = "low";

cyclonev_lcell_comb \Selector3~4 (
	.dataa(!at_sink_ready_s1),
	.datab(!\sink_state.run1~q ),
	.datac(!sink_valid),
	.datad(!\sink_state.stall~q ),
	.datae(!sink_sop),
	.dataf(!\sink_state.st_err~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~4 .extended_lut = "off";
defparam \Selector3~4 .lut_mask = 64'hFFFF7FDFFFFFFFFF;
defparam \Selector3~4 .shared_arith = "off";

cyclonev_lcell_comb \count~0 (
	.dataa(!\max_reached~q ),
	.datab(!\Selector3~6_combout ),
	.datac(!\count[0]~q ),
	.datad(!\Selector3~3_combout ),
	.datae(!\Selector3~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~0 .extended_lut = "off";
defparam \count~0 .lut_mask = 64'hFFFFFFB8FFFFFFB8;
defparam \count~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~1 (
	.dataa(!sink_error_0),
	.datab(!sink_error_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Selector2~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~6 (
	.dataa(!sink_valid),
	.datab(!\Selector2~1_combout ),
	.datac(!sink_sop),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~6 .extended_lut = "off";
defparam \Selector2~6 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Selector2~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~4 (
	.dataa(!\sink_state.run1~q ),
	.datab(!\sink_state.stall~q ),
	.datac(!at_sink_ready_s1),
	.datad(!\max_reached~q ),
	.datae(!sink_eop),
	.dataf(!\Selector2~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~4 .extended_lut = "off";
defparam \Selector2~4 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \Selector2~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~2 (
	.dataa(!at_sink_ready_s1),
	.datab(!\sink_state.run1~q ),
	.datac(!sink_valid),
	.datad(!\Selector2~1_combout ),
	.datae(!\sink_state.stall~q ),
	.dataf(!sink_sop),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'hFFFFDFFFFFFFFFFF;
defparam \Selector2~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~1 (
	.dataa(!sink_valid),
	.datab(!sink_error_0),
	.datac(!sink_error_1),
	.datad(!sink_sop),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Selector4~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!\max_reached~q ),
	.datab(!sink_eop),
	.datac(!at_sink_ready_s1),
	.datad(!\sink_state.run1~q ),
	.datae(!\sink_state.stall~q ),
	.dataf(!\Selector4~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \count[0]~1 (
	.dataa(!\Selector3~6_combout ),
	.datab(!\Selector2~4_combout ),
	.datac(!\Selector2~2_combout ),
	.datad(!\Selector3~3_combout ),
	.datae(!\Selector3~4_combout ),
	.dataf(!\Selector4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[0]~1 .extended_lut = "off";
defparam \count[0]~1 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \count[0]~1 .shared_arith = "off";

dffeas \count[0] (
	.clk(clk),
	.d(\count~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~1_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

cyclonev_lcell_comb \count~5 (
	.dataa(!\max_reached~q ),
	.datab(!\Selector3~6_combout ),
	.datac(!\count[1]~q ),
	.datad(!\count[0]~q ),
	.datae(!\Selector3~3_combout ),
	.dataf(!\Selector3~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~5 .extended_lut = "off";
defparam \count~5 .lut_mask = 64'hFFFFFFFFFFFFEBBE;
defparam \count~5 .shared_arith = "off";

dffeas \count[1] (
	.clk(clk),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~1_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \count~6 (
	.dataa(!\count[0]~q ),
	.datab(!\count[1]~q ),
	.datac(!\Selector3~3_combout ),
	.datad(!\count[2]~q ),
	.datae(!\Selector3~6_combout ),
	.dataf(!\max_reached~q ),
	.datag(!\Selector3~4_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~6 .extended_lut = "on";
defparam \count~6 .lut_mask = 64'h9F6F9F6F9F6F9F6F;
defparam \count~6 .shared_arith = "off";

dffeas \count[2] (
	.clk(clk),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~1_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\count[3]~q ),
	.datab(!\count[2]~q ),
	.datac(!\count[1]~q ),
	.datad(!\count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6996699669966996;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \count~4 (
	.dataa(!\max_reached~q ),
	.datab(!\Selector3~6_combout ),
	.datac(!\Selector3~3_combout ),
	.datad(!\Selector3~4_combout ),
	.datae(!\Add0~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~4 .extended_lut = "off";
defparam \count~4 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \count~4 .shared_arith = "off";

dffeas \count[3] (
	.clk(clk),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~1_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\count[4]~q ),
	.datab(!\count[3]~q ),
	.datac(!\count[2]~q ),
	.datad(!\count[1]~q ),
	.datae(!\count[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h9669699696696996;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \count~3 (
	.dataa(!\max_reached~q ),
	.datab(!\Selector3~6_combout ),
	.datac(!\Selector3~3_combout ),
	.datad(!\Selector3~4_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~3 .extended_lut = "off";
defparam \count~3 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \count~3 .shared_arith = "off";

dffeas \count[4] (
	.clk(clk),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~1_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\count[4]~q ),
	.datab(!\count[3]~q ),
	.datac(!\count[2]~q ),
	.datad(!\count[1]~q ),
	.datae(!\count[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \count~2 (
	.dataa(!\max_reached~q ),
	.datab(!\Selector3~6_combout ),
	.datac(!\count[5]~q ),
	.datad(!\Selector3~3_combout ),
	.datae(!\Selector3~4_combout ),
	.dataf(!\Add0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count~2 .extended_lut = "off";
defparam \count~2 .lut_mask = 64'hFFFFFFEBFFFFFFBE;
defparam \count~2 .shared_arith = "off";

dffeas \count[5] (
	.clk(clk),
	.d(\count~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~1_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

cyclonev_lcell_comb \max_reached~0 (
	.dataa(!\count[5]~q ),
	.datab(!\count[4]~q ),
	.datac(!\count[3]~q ),
	.datad(!\count[2]~q ),
	.datae(!\count[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\max_reached~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \max_reached~0 .extended_lut = "off";
defparam \max_reached~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \max_reached~0 .shared_arith = "off";

cyclonev_lcell_comb \max_reached~1 (
	.dataa(!\max_reached~q ),
	.datab(!\Selector2~3_combout ),
	.datac(!\count[0]~q ),
	.datad(!\Selector3~5_combout ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\max_reached~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\max_reached~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \max_reached~1 .extended_lut = "off";
defparam \max_reached~1 .lut_mask = 64'hFDF7F7FDFFFFFFFF;
defparam \max_reached~1 .shared_arith = "off";

dffeas max_reached(
	.clk(clk),
	.d(\max_reached~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\max_reached~q ),
	.prn(vcc));
defparam max_reached.is_wysiwyg = "true";
defparam max_reached.power_up = "low";

cyclonev_lcell_comb \Selector2~5 (
	.dataa(!sink_eop),
	.datab(!sink_valid),
	.datac(!\Selector2~1_combout ),
	.datad(!sink_sop),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~5 .extended_lut = "off";
defparam \Selector2~5 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Selector2~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~3 (
	.dataa(!at_sink_ready_s1),
	.datab(!\max_reached~q ),
	.datac(!\sink_state.stall~q ),
	.datad(!\sink_state.run1~q ),
	.datae(!sink_sop),
	.dataf(!\Selector2~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~3 .extended_lut = "off";
defparam \Selector2~3 .lut_mask = 64'hFDDFDFFDFFFFFFFF;
defparam \Selector2~3 .shared_arith = "off";

dffeas \sink_state.run1 (
	.clk(clk),
	.d(\Selector2~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.run1~q ),
	.prn(vcc));
defparam \sink_state.run1 .is_wysiwyg = "true";
defparam \sink_state.run1 .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\sink_state.run1~q ),
	.datab(!\sink_state.stall~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\sink_comb_update_2~0_combout ),
	.datab(!\Selector2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Selector1~0 .shared_arith = "off";

dffeas \sink_state.stall (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.stall~q ),
	.prn(vcc));
defparam \sink_state.stall .is_wysiwyg = "true";
defparam \sink_state.stall .power_up = "low";

cyclonev_lcell_comb \packet_error_int~0 (
	.dataa(!\max_reached~q ),
	.datab(!sink_eop),
	.datac(!sink_valid),
	.datad(!at_sink_ready_s1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_error_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_error_int~0 .extended_lut = "off";
defparam \packet_error_int~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \packet_error_int~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!at_sink_ready_s1),
	.datab(!\sink_state.run1~q ),
	.datac(!\max_reached~q ),
	.datad(!sink_eop),
	.datae(!sink_valid),
	.dataf(!sink_sop),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'hFFFFFFFF7FF7FFFF;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!sink_error_1),
	.datab(!\at_sink_error_int~0_combout ),
	.datac(!\sink_state.stall~q ),
	.datad(!sink_sop),
	.datae(!\packet_error_int~0_combout ),
	.dataf(!\Selector5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'hDF1FFFFFFFFFFFFF;
defparam \Selector5~1 .shared_arith = "off";

dffeas \sink_state.end1 (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.end1~q ),
	.prn(vcc));
defparam \sink_state.end1 .is_wysiwyg = "true";
defparam \sink_state.end1 .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\sink_state.end1~q ),
	.datab(!\sink_comb_update_2~0_combout ),
	.datac(!\sink_state.start~q ),
	.datad(!\sink_state.st_err~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \Selector0~0 .shared_arith = "off";

dffeas \sink_state.start (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_state.start~q ),
	.prn(vcc));
defparam \sink_state.start .is_wysiwyg = "true";
defparam \sink_state.start .power_up = "low";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!at_sink_ready_s1),
	.datab(!\sink_state.end1~q ),
	.datac(!sink_valid),
	.datad(!sink_sop),
	.datae(!\sink_state.start~q ),
	.dataf(!\sink_state.st_err~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \Selector6~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~1 (
	.dataa(!at_sink_ready_s1),
	.datab(!\max_reached~q ),
	.datac(!sink_eop),
	.datad(!sink_valid),
	.datae(!sink_sop),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \Selector6~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~2 (
	.dataa(!sink_error_0),
	.datab(!\at_sink_error_int~0_combout ),
	.datac(!\Selector2~0_combout ),
	.datad(!\Selector6~0_combout ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~2 .extended_lut = "off";
defparam \Selector6~2 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \Selector6~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!\out_cnt[5]~q ),
	.datab(!\out_cnt[4]~q ),
	.datac(!\out_cnt[3]~q ),
	.datad(!\out_cnt[2]~q ),
	.datae(!\out_cnt[1]~q ),
	.dataf(!\out_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal1~0 .shared_arith = "off";

endmodule

module IFFT_scfifo_1 (
	q,
	dffe_af,
	counter_reg_bit_0,
	empty_dff,
	sink_out_stateempty_and_ready,
	Selector7,
	sink_stall,
	Selector71,
	wrreq,
	Selector72,
	out_cnt_0,
	rdreq,
	data,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q;
output 	dffe_af;
output 	counter_reg_bit_0;
output 	empty_dff;
input 	sink_out_stateempty_and_ready;
input 	Selector7;
input 	sink_stall;
input 	Selector71;
input 	wrreq;
input 	Selector72;
input 	out_cnt_0;
input 	rdreq;
input 	[17:0] data;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IFFT_scfifo_d9p1 auto_generated(
	.q({q_unconnected_wire_17,q_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.dffe_af1(dffe_af),
	.counter_reg_bit_0(counter_reg_bit_0),
	.empty_dff(empty_dff),
	.sink_out_stateempty_and_ready(sink_out_stateempty_and_ready),
	.Selector7(Selector7),
	.sink_stall(sink_stall),
	.Selector71(Selector71),
	.wrreq(wrreq),
	.Selector72(Selector72),
	.out_cnt_0(out_cnt_0),
	.rdreq(rdreq),
	.data({gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module IFFT_scfifo_d9p1 (
	q,
	dffe_af1,
	counter_reg_bit_0,
	empty_dff,
	sink_out_stateempty_and_ready,
	Selector7,
	sink_stall,
	Selector71,
	wrreq,
	Selector72,
	out_cnt_0,
	rdreq,
	data,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q;
output 	dffe_af1;
output 	counter_reg_bit_0;
output 	empty_dff;
input 	sink_out_stateempty_and_ready;
input 	Selector7;
input 	sink_stall;
input 	Selector71;
input 	wrreq;
input 	Selector72;
input 	out_cnt_0;
input 	rdreq;
input 	[17:0] data;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;


IFFT_a_dpfifo_1je1 dpfifo(
	.q({q_unconnected_wire_17,q_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.counter_reg_bit_0(counter_reg_bit_0),
	.empty_dff1(empty_dff),
	.sink_out_stateempty_and_ready(sink_out_stateempty_and_ready),
	.Selector7(Selector7),
	.sink_stall(sink_stall),
	.Selector71(Selector71),
	.wreq(wrreq),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.Selector72(Selector72),
	.out_cnt_0(out_cnt_0),
	.rreq(rdreq),
	.data({gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock),
	.reset_n(reset_n));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

cyclonev_lcell_comb \dffe_af~0 (
	.dataa(!\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(!\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~0 .extended_lut = "off";
defparam \dffe_af~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \dffe_af~0 .shared_arith = "off";

cyclonev_lcell_comb \dffe_af~1 (
	.dataa(!dffe_af1),
	.datab(!counter_reg_bit_0),
	.datac(!Selector7),
	.datad(!Selector71),
	.datae(!wrreq),
	.dataf(!\dffe_af~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~1 .extended_lut = "off";
defparam \dffe_af~1 .lut_mask = 64'hFFFFFFDDFFFFFFF5;
defparam \dffe_af~1 .shared_arith = "off";

endmodule

module IFFT_a_dpfifo_1je1 (
	q,
	counter_reg_bit_0,
	empty_dff1,
	sink_out_stateempty_and_ready,
	Selector7,
	sink_stall,
	Selector71,
	wreq,
	counter_reg_bit_2,
	counter_reg_bit_1,
	Selector72,
	out_cnt_0,
	rreq,
	data,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q;
output 	counter_reg_bit_0;
output 	empty_dff1;
input 	sink_out_stateempty_and_ready;
input 	Selector7;
input 	sink_stall;
input 	Selector71;
input 	wreq;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	Selector72;
input 	out_cnt_0;
input 	rreq;
input 	[17:0] data;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \low_addressa[0]~q ;
wire \ram_read_address[0]~0_combout ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \_~4_combout ;
wire \_~3_combout ;
wire \usedw_is_0_dff~q ;
wire \_~1_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_is_1_dff~q ;
wire \_~2_combout ;


IFFT_altsyncram_afp1 FIFOram(
	.q_b({q_b_unconnected_wire_17,q_b_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren_a(wreq),
	.clocken1(rreq),
	.data_a({gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

IFFT_cntr_ggb wr_ptr(
	.fifo_wrreq(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.clock(clock),
	.reset_n(reset_n));

IFFT_cntr_sg7 usedw_counter(
	.counter_reg_bit_0(counter_reg_bit_0),
	.fifo_wrreq(wreq),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	._(\_~0_combout ),
	.clock(clock),
	.reset_n(reset_n));

IFFT_cntr_fgb rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	._(\_~4_combout ),
	.clock(clock),
	.reset_n(reset_n));

cyclonev_lcell_comb \_~0 (
	.dataa(!sink_stall),
	.datab(!sink_out_stateempty_and_ready),
	.datac(!Selector72),
	.datad(!wreq),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h6996699669966996;
defparam \_~0 .shared_arith = "off";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\ram_read_address[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

cyclonev_lcell_comb \ram_read_address[0]~0 (
	.dataa(!sink_stall),
	.datab(!sink_out_stateempty_and_ready),
	.datac(!Selector72),
	.datad(!out_cnt_0),
	.datae(!\low_addressa[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[0]~0 .extended_lut = "off";
defparam \ram_read_address[0]~0 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \ram_read_address[0]~0 .shared_arith = "off";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\ram_read_address[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cyclonev_lcell_comb \ram_read_address[1]~1 (
	.dataa(!sink_stall),
	.datab(!sink_out_stateempty_and_ready),
	.datac(!Selector72),
	.datad(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datae(!\low_addressa[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[1]~1 .extended_lut = "off";
defparam \ram_read_address[1]~1 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[1]~1 .shared_arith = "off";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\ram_read_address[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cyclonev_lcell_comb \ram_read_address[2]~2 (
	.dataa(!sink_stall),
	.datab(!sink_out_stateempty_and_ready),
	.datac(!Selector72),
	.datad(!\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datae(!\low_addressa[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[2]~2 .extended_lut = "off";
defparam \ram_read_address[2]~2 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \ram_read_address[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \_~4 (
	.dataa(!sink_stall),
	.datab(!sink_out_stateempty_and_ready),
	.datac(!Selector72),
	.datad(!out_cnt_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~4 .extended_lut = "off";
defparam \_~4 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \_~4 .shared_arith = "off";

dffeas empty_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cyclonev_lcell_comb \_~3 (
	.dataa(!sink_stall),
	.datab(!sink_out_stateempty_and_ready),
	.datac(!Selector72),
	.datad(!wreq),
	.datae(!\usedw_is_1_dff~q ),
	.dataf(!\usedw_is_0_dff~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~3 .extended_lut = "off";
defparam \_~3 .lut_mask = 64'hFFFF6996FFFFFFFF;
defparam \_~3 .shared_arith = "off";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\_~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter_reg_bit_0),
	.datab(!counter_reg_bit_2),
	.datac(!counter_reg_bit_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \usedw_will_be_1~0 (
	.dataa(!Selector7),
	.datab(!Selector71),
	.datac(!wreq),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(!\_~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \usedw_will_be_1~0 .extended_lut = "off";
defparam \usedw_will_be_1~0 .lut_mask = 64'hFFFF96FFFFFFFFFF;
defparam \usedw_will_be_1~0 .shared_arith = "off";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cyclonev_lcell_comb \_~2 (
	.dataa(!Selector7),
	.datab(!Selector71),
	.datac(!wreq),
	.datad(!\usedw_is_1_dff~q ),
	.datae(!\usedw_is_0_dff~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \_~2 .shared_arith = "off";

endmodule

module IFFT_altsyncram_afp1 (
	q_b,
	wren_a,
	clocken1,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[17:0] q_b;
input 	wren_a;
input 	clocken1;
input 	[17:0] data_a;
input 	[2:0] address_a;
input 	[2:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 18;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 18;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 18;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 18;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 18;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 18;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 18;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 18;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 18;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 18;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 18;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 18;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 18;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 18;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 18;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 18;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 18;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 18;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 18;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 18;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 18;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 18;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 18;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 18;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 18;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 18;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 18;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 18;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 18;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 18;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IFFT_fft_ii_0:fft_ii_0|asj_fft_sglstream:asj_fft_sglstream_inst|auk_dspip_avalon_streaming_sink:auk_dsp_atlantic_sink_1|scfifo:\\normal_fifo:fifo_eab_on:in_fifo|scfifo_d9p1:auto_generated|a_dpfifo_1je1:dpfifo|altsyncram_afp1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 18;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 18;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module IFFT_cntr_fgb (
	counter_reg_bit_0,
	counter_reg_bit_1,
	_,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	_;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

endmodule

module IFFT_cntr_ggb (
	fifo_wrreq,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	fifo_wrreq;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!fifo_wrreq),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!fifo_wrreq),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!fifo_wrreq),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

endmodule

module IFFT_cntr_sg7 (
	counter_reg_bit_0,
	fifo_wrreq,
	counter_reg_bit_2,
	counter_reg_bit_1,
	_,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
input 	fifo_wrreq;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	_;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!fifo_wrreq),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h0000FF00000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!fifo_wrreq),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h0000FF00000000FF;
defparam counter_comb_bita2.shared_arith = "off";

endmodule

module IFFT_auk_dspip_avalon_streaming_source (
	at_source_data_14,
	at_source_data_15,
	at_source_data_16,
	at_source_data_17,
	at_source_data_18,
	at_source_data_19,
	at_source_data_20,
	at_source_data_21,
	at_source_data_6,
	at_source_data_7,
	at_source_data_8,
	at_source_data_9,
	at_source_data_10,
	at_source_data_11,
	at_source_data_12,
	at_source_data_13,
	at_source_data_0,
	at_source_data_1,
	at_source_data_2,
	at_source_data_3,
	at_source_data_4,
	at_source_data_5,
	master_source_ena,
	data,
	at_source_valid_s1,
	at_source_error_0,
	at_source_error_1,
	at_source_sop_s1,
	at_source_eop_s1,
	source_packet_error_1,
	source_packet_error_0,
	sink_stall_reg,
	source_stall_reg,
	sink_ready_ctrl_d,
	send_sop_s,
	sop,
	stall_controller_comb,
	data_count,
	source_stall_int_d1,
	stall_reg,
	Mux0,
	Mux01,
	Mux02,
	stall_controller_comb1,
	clk,
	reset_n,
	source_ready)/* synthesis synthesis_greybox=1 */;
output 	at_source_data_14;
output 	at_source_data_15;
output 	at_source_data_16;
output 	at_source_data_17;
output 	at_source_data_18;
output 	at_source_data_19;
output 	at_source_data_20;
output 	at_source_data_21;
output 	at_source_data_6;
output 	at_source_data_7;
output 	at_source_data_8;
output 	at_source_data_9;
output 	at_source_data_10;
output 	at_source_data_11;
output 	at_source_data_12;
output 	at_source_data_13;
output 	at_source_data_0;
output 	at_source_data_1;
output 	at_source_data_2;
output 	at_source_data_3;
output 	at_source_data_4;
output 	at_source_data_5;
input 	master_source_ena;
input 	[21:0] data;
output 	at_source_valid_s1;
output 	at_source_error_0;
output 	at_source_error_1;
output 	at_source_sop_s1;
output 	at_source_eop_s1;
input 	source_packet_error_1;
input 	source_packet_error_0;
input 	sink_stall_reg;
input 	source_stall_reg;
input 	sink_ready_ctrl_d;
input 	send_sop_s;
input 	sop;
output 	stall_controller_comb;
input 	[5:0] data_count;
output 	source_stall_int_d1;
input 	stall_reg;
output 	Mux0;
output 	Mux01;
output 	Mux02;
output 	stall_controller_comb1;
input 	clk;
input 	reset_n;
input 	source_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \packet_error0~combout ;
wire \valid_ctrl_inter1~0_combout ;
wire \Mux3~0_combout ;
wire \valid_ctrl_inter1~1_combout ;
wire \valid_ctrl_int1~q ;
wire \first_data~0_combout ;
wire \first_data~q ;
wire \valid_ctrl_inter~0_combout ;
wire \valid_ctrl_inter~1_combout ;
wire \valid_ctrl_int~q ;
wire \Mux2~3_combout ;
wire \was_stalled~0_combout ;
wire \was_stalled~1_combout ;
wire \was_stalled~q ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \data_int[14]~q ;
wire \Mux3~1_combout ;
wire \data_int1[14]~q ;
wire \data_select~0_combout ;
wire \Mux1~0_combout ;
wire \data_int[15]~q ;
wire \data_int1[15]~q ;
wire \data_int[16]~q ;
wire \data_int1[16]~q ;
wire \data_int[17]~q ;
wire \data_int1[17]~q ;
wire \data_int[18]~q ;
wire \data_int1[18]~q ;
wire \data_int[19]~q ;
wire \data_int1[19]~q ;
wire \data_int[20]~q ;
wire \data_int1[20]~q ;
wire \data_int[21]~q ;
wire \data_int1[21]~q ;
wire \data_int[6]~q ;
wire \data_int1[6]~q ;
wire \data_int[7]~q ;
wire \data_int1[7]~q ;
wire \data_int[8]~q ;
wire \data_int1[8]~q ;
wire \data_int[9]~q ;
wire \data_int1[9]~q ;
wire \data_int[10]~q ;
wire \data_int1[10]~q ;
wire \data_int[11]~q ;
wire \data_int1[11]~q ;
wire \data_int[12]~q ;
wire \data_int1[12]~q ;
wire \data_int[13]~q ;
wire \data_int1[13]~q ;
wire \data_int[0]~q ;
wire \data_int1[0]~q ;
wire \data_int[1]~q ;
wire \data_int1[1]~q ;
wire \data_int[2]~q ;
wire \data_int1[2]~q ;
wire \data_int[3]~q ;
wire \data_int1[3]~q ;
wire \data_int[4]~q ;
wire \data_int1[4]~q ;
wire \data_int[5]~q ;
wire \data_int1[5]~q ;
wire \at_source_valid_int~0_combout ;
wire \Selector1~1_combout ;
wire \data_count_int1[4]~q ;
wire \data_count_int[4]~q ;
wire \packet_multi:count_finished~0_combout ;
wire \data_count_int[3]~q ;
wire \data_count_int[2]~q ;
wire \data_count_int[1]~q ;
wire \data_count_int[0]~q ;
wire \data_count_int[5]~q ;
wire \packet_multi:count_finished~1_combout ;
wire \data_count_int1[3]~q ;
wire \data_count_int1[2]~q ;
wire \data_count_int1[1]~q ;
wire \data_count_int1[0]~q ;
wire \data_count_int1[5]~q ;
wire \packet_multi:count_finished~2_combout ;
wire \packet_multi:count_finished~combout ;
wire \source_comb_update_2~0_combout ;
wire \source_comb_update_2~2_combout ;
wire \source_comb_update_2~3_combout ;
wire \source_comb_update_2~1_combout ;
wire \packet_multi:source_state.run1~q ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \packet_multi:source_state.end1~q ;
wire \Selector0~0_combout ;
wire \packet_multi:source_state.st_err~q ;
wire \Selector0~1_combout ;
wire \packet_multi:source_state.start~q ;
wire \Selector1~3_combout ;
wire \Selector1~4_combout ;
wire \packet_multi:source_state.sop~q ;
wire \Selector2~0_combout ;
wire \Selector1~0_combout ;
wire \Selector1~2_combout ;
wire \at_source_valid_int~1_combout ;
wire \at_source_valid_int~2_combout ;
wire \at_source_valid_int~3_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;


dffeas \at_source_data[14] (
	.clk(clk),
	.d(\data_int[14]~q ),
	.asdata(\data_int1[14]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_14),
	.prn(vcc));
defparam \at_source_data[14] .is_wysiwyg = "true";
defparam \at_source_data[14] .power_up = "low";

dffeas \at_source_data[15] (
	.clk(clk),
	.d(\data_int[15]~q ),
	.asdata(\data_int1[15]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_15),
	.prn(vcc));
defparam \at_source_data[15] .is_wysiwyg = "true";
defparam \at_source_data[15] .power_up = "low";

dffeas \at_source_data[16] (
	.clk(clk),
	.d(\data_int[16]~q ),
	.asdata(\data_int1[16]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_16),
	.prn(vcc));
defparam \at_source_data[16] .is_wysiwyg = "true";
defparam \at_source_data[16] .power_up = "low";

dffeas \at_source_data[17] (
	.clk(clk),
	.d(\data_int[17]~q ),
	.asdata(\data_int1[17]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_17),
	.prn(vcc));
defparam \at_source_data[17] .is_wysiwyg = "true";
defparam \at_source_data[17] .power_up = "low";

dffeas \at_source_data[18] (
	.clk(clk),
	.d(\data_int[18]~q ),
	.asdata(\data_int1[18]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_18),
	.prn(vcc));
defparam \at_source_data[18] .is_wysiwyg = "true";
defparam \at_source_data[18] .power_up = "low";

dffeas \at_source_data[19] (
	.clk(clk),
	.d(\data_int[19]~q ),
	.asdata(\data_int1[19]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_19),
	.prn(vcc));
defparam \at_source_data[19] .is_wysiwyg = "true";
defparam \at_source_data[19] .power_up = "low";

dffeas \at_source_data[20] (
	.clk(clk),
	.d(\data_int[20]~q ),
	.asdata(\data_int1[20]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_20),
	.prn(vcc));
defparam \at_source_data[20] .is_wysiwyg = "true";
defparam \at_source_data[20] .power_up = "low";

dffeas \at_source_data[21] (
	.clk(clk),
	.d(\data_int[21]~q ),
	.asdata(\data_int1[21]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_21),
	.prn(vcc));
defparam \at_source_data[21] .is_wysiwyg = "true";
defparam \at_source_data[21] .power_up = "low";

dffeas \at_source_data[6] (
	.clk(clk),
	.d(\data_int[6]~q ),
	.asdata(\data_int1[6]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_6),
	.prn(vcc));
defparam \at_source_data[6] .is_wysiwyg = "true";
defparam \at_source_data[6] .power_up = "low";

dffeas \at_source_data[7] (
	.clk(clk),
	.d(\data_int[7]~q ),
	.asdata(\data_int1[7]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_7),
	.prn(vcc));
defparam \at_source_data[7] .is_wysiwyg = "true";
defparam \at_source_data[7] .power_up = "low";

dffeas \at_source_data[8] (
	.clk(clk),
	.d(\data_int[8]~q ),
	.asdata(\data_int1[8]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_8),
	.prn(vcc));
defparam \at_source_data[8] .is_wysiwyg = "true";
defparam \at_source_data[8] .power_up = "low";

dffeas \at_source_data[9] (
	.clk(clk),
	.d(\data_int[9]~q ),
	.asdata(\data_int1[9]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_9),
	.prn(vcc));
defparam \at_source_data[9] .is_wysiwyg = "true";
defparam \at_source_data[9] .power_up = "low";

dffeas \at_source_data[10] (
	.clk(clk),
	.d(\data_int[10]~q ),
	.asdata(\data_int1[10]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_10),
	.prn(vcc));
defparam \at_source_data[10] .is_wysiwyg = "true";
defparam \at_source_data[10] .power_up = "low";

dffeas \at_source_data[11] (
	.clk(clk),
	.d(\data_int[11]~q ),
	.asdata(\data_int1[11]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_11),
	.prn(vcc));
defparam \at_source_data[11] .is_wysiwyg = "true";
defparam \at_source_data[11] .power_up = "low";

dffeas \at_source_data[12] (
	.clk(clk),
	.d(\data_int[12]~q ),
	.asdata(\data_int1[12]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_12),
	.prn(vcc));
defparam \at_source_data[12] .is_wysiwyg = "true";
defparam \at_source_data[12] .power_up = "low";

dffeas \at_source_data[13] (
	.clk(clk),
	.d(\data_int[13]~q ),
	.asdata(\data_int1[13]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_13),
	.prn(vcc));
defparam \at_source_data[13] .is_wysiwyg = "true";
defparam \at_source_data[13] .power_up = "low";

dffeas \at_source_data[0] (
	.clk(clk),
	.d(\data_int[0]~q ),
	.asdata(\data_int1[0]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_0),
	.prn(vcc));
defparam \at_source_data[0] .is_wysiwyg = "true";
defparam \at_source_data[0] .power_up = "low";

dffeas \at_source_data[1] (
	.clk(clk),
	.d(\data_int[1]~q ),
	.asdata(\data_int1[1]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_1),
	.prn(vcc));
defparam \at_source_data[1] .is_wysiwyg = "true";
defparam \at_source_data[1] .power_up = "low";

dffeas \at_source_data[2] (
	.clk(clk),
	.d(\data_int[2]~q ),
	.asdata(\data_int1[2]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_2),
	.prn(vcc));
defparam \at_source_data[2] .is_wysiwyg = "true";
defparam \at_source_data[2] .power_up = "low";

dffeas \at_source_data[3] (
	.clk(clk),
	.d(\data_int[3]~q ),
	.asdata(\data_int1[3]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_3),
	.prn(vcc));
defparam \at_source_data[3] .is_wysiwyg = "true";
defparam \at_source_data[3] .power_up = "low";

dffeas \at_source_data[4] (
	.clk(clk),
	.d(\data_int[4]~q ),
	.asdata(\data_int1[4]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_4),
	.prn(vcc));
defparam \at_source_data[4] .is_wysiwyg = "true";
defparam \at_source_data[4] .power_up = "low";

dffeas \at_source_data[5] (
	.clk(clk),
	.d(\data_int[5]~q ),
	.asdata(\data_int1[5]~q ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\data_select~0_combout ),
	.ena(\Mux1~0_combout ),
	.q(at_source_data_5),
	.prn(vcc));
defparam \at_source_data[5] .is_wysiwyg = "true";
defparam \at_source_data[5] .power_up = "low";

dffeas at_source_valid_s(
	.clk(clk),
	.d(\at_source_valid_int~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_valid_s1),
	.prn(vcc));
defparam at_source_valid_s.is_wysiwyg = "true";
defparam at_source_valid_s.power_up = "low";

dffeas \at_source_error[0] (
	.clk(clk),
	.d(source_packet_error_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_0),
	.prn(vcc));
defparam \at_source_error[0] .is_wysiwyg = "true";
defparam \at_source_error[0] .power_up = "low";

dffeas \at_source_error[1] (
	.clk(clk),
	.d(source_packet_error_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_error_1),
	.prn(vcc));
defparam \at_source_error[1] .is_wysiwyg = "true";
defparam \at_source_error[1] .power_up = "low";

dffeas at_source_sop_s(
	.clk(clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_sop_s1),
	.prn(vcc));
defparam at_source_sop_s.is_wysiwyg = "true";
defparam at_source_sop_s.power_up = "low";

dffeas at_source_eop_s(
	.clk(clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(at_source_eop_s1),
	.prn(vcc));
defparam at_source_eop_s.is_wysiwyg = "true";
defparam at_source_eop_s.power_up = "low";

cyclonev_lcell_comb \stall_controller_comb~0 (
	.dataa(!sink_stall_reg),
	.datab(!source_stall_reg),
	.datac(!sink_ready_ctrl_d),
	.datad(!send_sop_s),
	.datae(!sop),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(stall_controller_comb),
	.sumout(),
	.cout(),
	.shareout());
defparam \stall_controller_comb~0 .extended_lut = "off";
defparam \stall_controller_comb~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \stall_controller_comb~0 .shared_arith = "off";

dffeas source_stall_int_d(
	.clk(clk),
	.d(Mux02),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_int_d1),
	.prn(vcc));
defparam source_stall_int_d.is_wysiwyg = "true";
defparam source_stall_int_d.power_up = "low";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\valid_ctrl_int~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~1 (
	.dataa(!source_ready),
	.datab(!\valid_ctrl_int~q ),
	.datac(!\first_data~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux01),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~1 .extended_lut = "off";
defparam \Mux0~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \Mux0~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~2 (
	.dataa(!at_source_valid_s1),
	.datab(!\was_stalled~q ),
	.datac(!master_source_ena),
	.datad(!stall_controller_comb),
	.datae(!Mux0),
	.dataf(!Mux01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux02),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~2 .extended_lut = "off";
defparam \Mux0~2 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \Mux0~2 .shared_arith = "off";

cyclonev_lcell_comb \stall_controller_comb~1 (
	.dataa(!\was_stalled~q ),
	.datab(!master_source_ena),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(stall_controller_comb1),
	.sumout(),
	.cout(),
	.shareout());
defparam \stall_controller_comb~1 .extended_lut = "off";
defparam \stall_controller_comb~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \stall_controller_comb~1 .shared_arith = "off";

cyclonev_lcell_comb packet_error0(
	.dataa(!source_packet_error_1),
	.datab(!source_packet_error_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_error0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam packet_error0.extended_lut = "off";
defparam packet_error0.lut_mask = 64'h7777777777777777;
defparam packet_error0.shared_arith = "off";

cyclonev_lcell_comb \valid_ctrl_inter1~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(gnd),
	.datad(!\first_data~q ),
	.datae(!\valid_ctrl_int1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_ctrl_inter1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_ctrl_inter1~0 .extended_lut = "off";
defparam \valid_ctrl_inter1~0 .lut_mask = 64'hFFEEFFFFFFEEFFFF;
defparam \valid_ctrl_inter1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\valid_ctrl_int~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \valid_ctrl_inter1~1 (
	.dataa(!\was_stalled~q ),
	.datab(!master_source_ena),
	.datac(!stall_controller_comb),
	.datad(!\valid_ctrl_inter1~0_combout ),
	.datae(!\Mux3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_ctrl_inter1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_ctrl_inter1~1 .extended_lut = "off";
defparam \valid_ctrl_inter1~1 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \valid_ctrl_inter1~1 .shared_arith = "off";

dffeas valid_ctrl_int1(
	.clk(clk),
	.d(\valid_ctrl_inter1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int1~q ),
	.prn(vcc));
defparam valid_ctrl_int1.is_wysiwyg = "true";
defparam valid_ctrl_int1.power_up = "low";

cyclonev_lcell_comb \first_data~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\first_data~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\first_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \first_data~0 .extended_lut = "off";
defparam \first_data~0 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \first_data~0 .shared_arith = "off";

dffeas first_data(
	.clk(clk),
	.d(\first_data~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\first_data~q ),
	.prn(vcc));
defparam first_data.is_wysiwyg = "true";
defparam first_data.power_up = "low";

cyclonev_lcell_comb \valid_ctrl_inter~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\packet_error0~combout ),
	.datac(!source_ready),
	.datad(!\valid_ctrl_int~q ),
	.datae(!\first_data~q ),
	.dataf(!\valid_ctrl_int1~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_ctrl_inter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_ctrl_inter~0 .extended_lut = "off";
defparam \valid_ctrl_inter~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \valid_ctrl_inter~0 .shared_arith = "off";

cyclonev_lcell_comb \valid_ctrl_inter~1 (
	.dataa(!\was_stalled~q ),
	.datab(!master_source_ena),
	.datac(!\Mux2~3_combout ),
	.datad(!stall_controller_comb),
	.datae(gnd),
	.dataf(!\valid_ctrl_inter~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\valid_ctrl_inter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \valid_ctrl_inter~1 .extended_lut = "off";
defparam \valid_ctrl_inter~1 .lut_mask = 64'hFFFBFFFBFFFFFFFF;
defparam \valid_ctrl_inter~1 .shared_arith = "off";

dffeas valid_ctrl_int(
	.clk(clk),
	.d(\valid_ctrl_inter~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\valid_ctrl_int~q ),
	.prn(vcc));
defparam valid_ctrl_int.is_wysiwyg = "true";
defparam valid_ctrl_int.power_up = "low";

cyclonev_lcell_comb \Mux2~3 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\valid_ctrl_int~q ),
	.datad(!\first_data~q ),
	.datae(!\valid_ctrl_int1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~3 .extended_lut = "off";
defparam \Mux2~3 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \Mux2~3 .shared_arith = "off";

cyclonev_lcell_comb \was_stalled~0 (
	.dataa(!sink_ready_ctrl_d),
	.datab(!send_sop_s),
	.datac(!sop),
	.datad(!source_stall_int_d1),
	.datae(!stall_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\was_stalled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \was_stalled~0 .extended_lut = "off";
defparam \was_stalled~0 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \was_stalled~0 .shared_arith = "off";

cyclonev_lcell_comb \was_stalled~1 (
	.dataa(!\was_stalled~q ),
	.datab(!master_source_ena),
	.datac(!\Mux2~3_combout ),
	.datad(!stall_controller_comb),
	.datae(!\was_stalled~0_combout ),
	.dataf(!\Mux3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\was_stalled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \was_stalled~1 .extended_lut = "off";
defparam \was_stalled~1 .lut_mask = 64'hFFFFFFF7FFFFFFFF;
defparam \was_stalled~1 .shared_arith = "off";

dffeas was_stalled(
	.clk(clk),
	.d(\was_stalled~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\was_stalled~q ),
	.prn(vcc));
defparam was_stalled.is_wysiwyg = "true";
defparam was_stalled.power_up = "low";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\valid_ctrl_int~q ),
	.datac(!\valid_ctrl_int1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~1 (
	.dataa(!at_source_valid_s1),
	.datab(!\first_data~q ),
	.datac(!\valid_ctrl_int1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~1 .extended_lut = "off";
defparam \Mux2~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Mux2~1 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~2 (
	.dataa(!source_ready),
	.datab(!\was_stalled~q ),
	.datac(!master_source_ena),
	.datad(!\Mux2~0_combout ),
	.datae(!\Mux2~1_combout ),
	.dataf(!stall_controller_comb),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~2 .extended_lut = "off";
defparam \Mux2~2 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \Mux2~2 .shared_arith = "off";

dffeas \data_int[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[14]~q ),
	.prn(vcc));
defparam \data_int[14] .is_wysiwyg = "true";
defparam \data_int[14] .power_up = "low";

cyclonev_lcell_comb \Mux3~1 (
	.dataa(!source_ready),
	.datab(!\valid_ctrl_int1~q ),
	.datac(!\was_stalled~q ),
	.datad(!master_source_ena),
	.datae(!\Mux2~0_combout ),
	.dataf(!stall_controller_comb),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~1 .extended_lut = "off";
defparam \Mux3~1 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Mux3~1 .shared_arith = "off";

dffeas \data_int1[14] (
	.clk(clk),
	.d(data[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[14]~q ),
	.prn(vcc));
defparam \data_int1[14] .is_wysiwyg = "true";
defparam \data_int1[14] .power_up = "low";

cyclonev_lcell_comb \data_select~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\first_data~q ),
	.datac(!\valid_ctrl_int1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_select~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_select~0 .extended_lut = "off";
defparam \data_select~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \data_select~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\valid_ctrl_int~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \Mux1~0 .shared_arith = "off";

dffeas \data_int[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[15]~q ),
	.prn(vcc));
defparam \data_int[15] .is_wysiwyg = "true";
defparam \data_int[15] .power_up = "low";

dffeas \data_int1[15] (
	.clk(clk),
	.d(data[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[15]~q ),
	.prn(vcc));
defparam \data_int1[15] .is_wysiwyg = "true";
defparam \data_int1[15] .power_up = "low";

dffeas \data_int[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[16]~q ),
	.prn(vcc));
defparam \data_int[16] .is_wysiwyg = "true";
defparam \data_int[16] .power_up = "low";

dffeas \data_int1[16] (
	.clk(clk),
	.d(data[16]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[16]~q ),
	.prn(vcc));
defparam \data_int1[16] .is_wysiwyg = "true";
defparam \data_int1[16] .power_up = "low";

dffeas \data_int[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[17]~q ),
	.prn(vcc));
defparam \data_int[17] .is_wysiwyg = "true";
defparam \data_int[17] .power_up = "low";

dffeas \data_int1[17] (
	.clk(clk),
	.d(data[17]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[17]~q ),
	.prn(vcc));
defparam \data_int1[17] .is_wysiwyg = "true";
defparam \data_int1[17] .power_up = "low";

dffeas \data_int[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[18]~q ),
	.prn(vcc));
defparam \data_int[18] .is_wysiwyg = "true";
defparam \data_int[18] .power_up = "low";

dffeas \data_int1[18] (
	.clk(clk),
	.d(data[18]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[18]~q ),
	.prn(vcc));
defparam \data_int1[18] .is_wysiwyg = "true";
defparam \data_int1[18] .power_up = "low";

dffeas \data_int[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[19]~q ),
	.prn(vcc));
defparam \data_int[19] .is_wysiwyg = "true";
defparam \data_int[19] .power_up = "low";

dffeas \data_int1[19] (
	.clk(clk),
	.d(data[19]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[19]~q ),
	.prn(vcc));
defparam \data_int1[19] .is_wysiwyg = "true";
defparam \data_int1[19] .power_up = "low";

dffeas \data_int[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[20]~q ),
	.prn(vcc));
defparam \data_int[20] .is_wysiwyg = "true";
defparam \data_int[20] .power_up = "low";

dffeas \data_int1[20] (
	.clk(clk),
	.d(data[20]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[20]~q ),
	.prn(vcc));
defparam \data_int1[20] .is_wysiwyg = "true";
defparam \data_int1[20] .power_up = "low";

dffeas \data_int[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[21]~q ),
	.prn(vcc));
defparam \data_int[21] .is_wysiwyg = "true";
defparam \data_int[21] .power_up = "low";

dffeas \data_int1[21] (
	.clk(clk),
	.d(data[21]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[21]~q ),
	.prn(vcc));
defparam \data_int1[21] .is_wysiwyg = "true";
defparam \data_int1[21] .power_up = "low";

dffeas \data_int[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[6]~q ),
	.prn(vcc));
defparam \data_int[6] .is_wysiwyg = "true";
defparam \data_int[6] .power_up = "low";

dffeas \data_int1[6] (
	.clk(clk),
	.d(data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[6]~q ),
	.prn(vcc));
defparam \data_int1[6] .is_wysiwyg = "true";
defparam \data_int1[6] .power_up = "low";

dffeas \data_int[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[7]~q ),
	.prn(vcc));
defparam \data_int[7] .is_wysiwyg = "true";
defparam \data_int[7] .power_up = "low";

dffeas \data_int1[7] (
	.clk(clk),
	.d(data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[7]~q ),
	.prn(vcc));
defparam \data_int1[7] .is_wysiwyg = "true";
defparam \data_int1[7] .power_up = "low";

dffeas \data_int[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[8]~q ),
	.prn(vcc));
defparam \data_int[8] .is_wysiwyg = "true";
defparam \data_int[8] .power_up = "low";

dffeas \data_int1[8] (
	.clk(clk),
	.d(data[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[8]~q ),
	.prn(vcc));
defparam \data_int1[8] .is_wysiwyg = "true";
defparam \data_int1[8] .power_up = "low";

dffeas \data_int[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[9]~q ),
	.prn(vcc));
defparam \data_int[9] .is_wysiwyg = "true";
defparam \data_int[9] .power_up = "low";

dffeas \data_int1[9] (
	.clk(clk),
	.d(data[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[9]~q ),
	.prn(vcc));
defparam \data_int1[9] .is_wysiwyg = "true";
defparam \data_int1[9] .power_up = "low";

dffeas \data_int[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[10]~q ),
	.prn(vcc));
defparam \data_int[10] .is_wysiwyg = "true";
defparam \data_int[10] .power_up = "low";

dffeas \data_int1[10] (
	.clk(clk),
	.d(data[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[10]~q ),
	.prn(vcc));
defparam \data_int1[10] .is_wysiwyg = "true";
defparam \data_int1[10] .power_up = "low";

dffeas \data_int[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[11]~q ),
	.prn(vcc));
defparam \data_int[11] .is_wysiwyg = "true";
defparam \data_int[11] .power_up = "low";

dffeas \data_int1[11] (
	.clk(clk),
	.d(data[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[11]~q ),
	.prn(vcc));
defparam \data_int1[11] .is_wysiwyg = "true";
defparam \data_int1[11] .power_up = "low";

dffeas \data_int[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[12]~q ),
	.prn(vcc));
defparam \data_int[12] .is_wysiwyg = "true";
defparam \data_int[12] .power_up = "low";

dffeas \data_int1[12] (
	.clk(clk),
	.d(data[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[12]~q ),
	.prn(vcc));
defparam \data_int1[12] .is_wysiwyg = "true";
defparam \data_int1[12] .power_up = "low";

dffeas \data_int[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[13]~q ),
	.prn(vcc));
defparam \data_int[13] .is_wysiwyg = "true";
defparam \data_int[13] .power_up = "low";

dffeas \data_int1[13] (
	.clk(clk),
	.d(data[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[13]~q ),
	.prn(vcc));
defparam \data_int1[13] .is_wysiwyg = "true";
defparam \data_int1[13] .power_up = "low";

dffeas \data_int[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[0]~q ),
	.prn(vcc));
defparam \data_int[0] .is_wysiwyg = "true";
defparam \data_int[0] .power_up = "low";

dffeas \data_int1[0] (
	.clk(clk),
	.d(data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[0]~q ),
	.prn(vcc));
defparam \data_int1[0] .is_wysiwyg = "true";
defparam \data_int1[0] .power_up = "low";

dffeas \data_int[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[1]~q ),
	.prn(vcc));
defparam \data_int[1] .is_wysiwyg = "true";
defparam \data_int[1] .power_up = "low";

dffeas \data_int1[1] (
	.clk(clk),
	.d(data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[1]~q ),
	.prn(vcc));
defparam \data_int1[1] .is_wysiwyg = "true";
defparam \data_int1[1] .power_up = "low";

dffeas \data_int[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[2]~q ),
	.prn(vcc));
defparam \data_int[2] .is_wysiwyg = "true";
defparam \data_int[2] .power_up = "low";

dffeas \data_int1[2] (
	.clk(clk),
	.d(data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[2]~q ),
	.prn(vcc));
defparam \data_int1[2] .is_wysiwyg = "true";
defparam \data_int1[2] .power_up = "low";

dffeas \data_int[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[3]~q ),
	.prn(vcc));
defparam \data_int[3] .is_wysiwyg = "true";
defparam \data_int[3] .power_up = "low";

dffeas \data_int1[3] (
	.clk(clk),
	.d(data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[3]~q ),
	.prn(vcc));
defparam \data_int1[3] .is_wysiwyg = "true";
defparam \data_int1[3] .power_up = "low";

dffeas \data_int[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[4]~q ),
	.prn(vcc));
defparam \data_int[4] .is_wysiwyg = "true";
defparam \data_int[4] .power_up = "low";

dffeas \data_int1[4] (
	.clk(clk),
	.d(data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[4]~q ),
	.prn(vcc));
defparam \data_int1[4] .is_wysiwyg = "true";
defparam \data_int1[4] .power_up = "low";

dffeas \data_int[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_int[5]~q ),
	.prn(vcc));
defparam \data_int[5] .is_wysiwyg = "true";
defparam \data_int[5] .power_up = "low";

dffeas \data_int1[5] (
	.clk(clk),
	.d(data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_int1[5]~q ),
	.prn(vcc));
defparam \data_int1[5] .is_wysiwyg = "true";
defparam \data_int1[5] .power_up = "low";

cyclonev_lcell_comb \at_source_valid_int~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_packet_error_1),
	.datac(!source_packet_error_0),
	.datad(!source_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\at_source_valid_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \at_source_valid_int~0 .extended_lut = "off";
defparam \at_source_valid_int~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \at_source_valid_int~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!source_packet_error_1),
	.datab(!source_packet_error_0),
	.datac(!\packet_multi:source_state.sop~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Selector1~1 .shared_arith = "off";

dffeas \data_count_int1[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[4]~q ),
	.prn(vcc));
defparam \data_count_int1[4] .is_wysiwyg = "true";
defparam \data_count_int1[4] .power_up = "low";

dffeas \data_count_int[4] (
	.clk(clk),
	.d(data_count[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_count_int[4]~q ),
	.prn(vcc));
defparam \data_count_int[4] .is_wysiwyg = "true";
defparam \data_count_int[4] .power_up = "low";

cyclonev_lcell_comb \packet_multi:count_finished~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\valid_ctrl_int~q ),
	.datac(!\first_data~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(!\data_count_int1[4]~q ),
	.dataf(!\data_count_int[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_multi:count_finished~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_multi:count_finished~0 .extended_lut = "off";
defparam \packet_multi:count_finished~0 .lut_mask = 64'hB77BFFFFFFFFFFFF;
defparam \packet_multi:count_finished~0 .shared_arith = "off";

dffeas \data_count_int[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_count_int[3]~q ),
	.prn(vcc));
defparam \data_count_int[3] .is_wysiwyg = "true";
defparam \data_count_int[3] .power_up = "low";

dffeas \data_count_int[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_count_int[2]~q ),
	.prn(vcc));
defparam \data_count_int[2] .is_wysiwyg = "true";
defparam \data_count_int[2] .power_up = "low";

dffeas \data_count_int[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_count_int[1]~q ),
	.prn(vcc));
defparam \data_count_int[1] .is_wysiwyg = "true";
defparam \data_count_int[1] .power_up = "low";

dffeas \data_count_int[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_count_int[0]~q ),
	.prn(vcc));
defparam \data_count_int[0] .is_wysiwyg = "true";
defparam \data_count_int[0] .power_up = "low";

dffeas \data_count_int[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux2~2_combout ),
	.q(\data_count_int[5]~q ),
	.prn(vcc));
defparam \data_count_int[5] .is_wysiwyg = "true";
defparam \data_count_int[5] .power_up = "low";

cyclonev_lcell_comb \packet_multi:count_finished~1 (
	.dataa(!\data_count_int[3]~q ),
	.datab(!\data_count_int[2]~q ),
	.datac(!\data_count_int[1]~q ),
	.datad(!\data_count_int[0]~q ),
	.datae(!\data_count_int[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_multi:count_finished~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_multi:count_finished~1 .extended_lut = "off";
defparam \packet_multi:count_finished~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \packet_multi:count_finished~1 .shared_arith = "off";

dffeas \data_count_int1[3] (
	.clk(clk),
	.d(data_count[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[3]~q ),
	.prn(vcc));
defparam \data_count_int1[3] .is_wysiwyg = "true";
defparam \data_count_int1[3] .power_up = "low";

dffeas \data_count_int1[2] (
	.clk(clk),
	.d(data_count[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[2]~q ),
	.prn(vcc));
defparam \data_count_int1[2] .is_wysiwyg = "true";
defparam \data_count_int1[2] .power_up = "low";

dffeas \data_count_int1[1] (
	.clk(clk),
	.d(data_count[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[1]~q ),
	.prn(vcc));
defparam \data_count_int1[1] .is_wysiwyg = "true";
defparam \data_count_int1[1] .power_up = "low";

dffeas \data_count_int1[0] (
	.clk(clk),
	.d(data_count[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[0]~q ),
	.prn(vcc));
defparam \data_count_int1[0] .is_wysiwyg = "true";
defparam \data_count_int1[0] .power_up = "low";

dffeas \data_count_int1[5] (
	.clk(clk),
	.d(data_count[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux3~1_combout ),
	.q(\data_count_int1[5]~q ),
	.prn(vcc));
defparam \data_count_int1[5] .is_wysiwyg = "true";
defparam \data_count_int1[5] .power_up = "low";

cyclonev_lcell_comb \packet_multi:count_finished~2 (
	.dataa(!\data_count_int1[3]~q ),
	.datab(!\data_count_int1[2]~q ),
	.datac(!\data_count_int1[1]~q ),
	.datad(!\data_count_int1[0]~q ),
	.datae(!\data_count_int1[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_multi:count_finished~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_multi:count_finished~2 .extended_lut = "off";
defparam \packet_multi:count_finished~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \packet_multi:count_finished~2 .shared_arith = "off";

cyclonev_lcell_comb \packet_multi:count_finished (
	.dataa(!\packet_multi:count_finished~0_combout ),
	.datab(!at_source_valid_s1),
	.datac(!\first_data~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(!\packet_multi:count_finished~1_combout ),
	.dataf(!\packet_multi:count_finished~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_multi:count_finished~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_multi:count_finished .extended_lut = "off";
defparam \packet_multi:count_finished .lut_mask = 64'hD77DFFFFFFFFFFFF;
defparam \packet_multi:count_finished .shared_arith = "off";

cyclonev_lcell_comb \source_comb_update_2~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\valid_ctrl_int~q ),
	.datac(!\first_data~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(!\data_count_int1[4]~q ),
	.dataf(!\data_count_int[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_comb_update_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_comb_update_2~0 .extended_lut = "off";
defparam \source_comb_update_2~0 .lut_mask = 64'hFFFFFFFFFFFFB77B;
defparam \source_comb_update_2~0 .shared_arith = "off";

cyclonev_lcell_comb \source_comb_update_2~2 (
	.dataa(!\data_count_int[3]~q ),
	.datab(!\data_count_int[2]~q ),
	.datac(!\data_count_int[1]~q ),
	.datad(!\data_count_int[0]~q ),
	.datae(!\data_count_int[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_comb_update_2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_comb_update_2~2 .extended_lut = "off";
defparam \source_comb_update_2~2 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \source_comb_update_2~2 .shared_arith = "off";

cyclonev_lcell_comb \source_comb_update_2~3 (
	.dataa(!\data_count_int1[3]~q ),
	.datab(!\data_count_int1[2]~q ),
	.datac(!\data_count_int1[1]~q ),
	.datad(!\data_count_int1[0]~q ),
	.datae(!\data_count_int1[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_comb_update_2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_comb_update_2~3 .extended_lut = "off";
defparam \source_comb_update_2~3 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \source_comb_update_2~3 .shared_arith = "off";

cyclonev_lcell_comb \source_comb_update_2~1 (
	.dataa(!\source_comb_update_2~0_combout ),
	.datab(!at_source_valid_s1),
	.datac(!\first_data~q ),
	.datad(!\valid_ctrl_int1~q ),
	.datae(!\source_comb_update_2~2_combout ),
	.dataf(!\source_comb_update_2~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\source_comb_update_2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \source_comb_update_2~1 .extended_lut = "off";
defparam \source_comb_update_2~1 .lut_mask = 64'hD77DFFFFFFFFFFFF;
defparam \source_comb_update_2~1 .shared_arith = "off";

dffeas \packet_multi:source_state.run1 (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.run1~q ),
	.prn(vcc));
defparam \packet_multi:source_state.run1 .is_wysiwyg = "true";
defparam \packet_multi:source_state.run1 .power_up = "low";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\packet_multi:source_state.sop~q ),
	.datab(!\packet_multi:source_state.run1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!at_source_valid_s1),
	.datab(!\packet_error0~combout ),
	.datac(!source_ready),
	.datad(!\packet_multi:count_finished~combout ),
	.datae(!\packet_multi:source_state.end1~q ),
	.dataf(!\Selector3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'hFFFFFFFFACFFFFFF;
defparam \Selector3~1 .shared_arith = "off";

dffeas \packet_multi:source_state.end1 (
	.clk(clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.end1~q ),
	.prn(vcc));
defparam \packet_multi:source_state.end1 .is_wysiwyg = "true";
defparam \packet_multi:source_state.end1 .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\packet_multi:source_state.start~q ),
	.datad(!\packet_multi:source_state.end1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \Selector0~0 .shared_arith = "off";

dffeas \packet_multi:source_state.st_err (
	.clk(clk),
	.d(\packet_error0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.st_err~q ),
	.prn(vcc));
defparam \packet_multi:source_state.st_err .is_wysiwyg = "true";
defparam \packet_multi:source_state.st_err .power_up = "low";

cyclonev_lcell_comb \Selector0~1 (
	.dataa(!\packet_error0~combout ),
	.datab(!\Selector0~0_combout ),
	.datac(!\source_comb_update_2~1_combout ),
	.datad(!\packet_multi:source_state.st_err~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \Selector0~1 .shared_arith = "off";

dffeas \packet_multi:source_state.start (
	.clk(clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.start~q ),
	.prn(vcc));
defparam \packet_multi:source_state.start .is_wysiwyg = "true";
defparam \packet_multi:source_state.start .power_up = "low";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!at_source_valid_s1),
	.datab(!source_packet_error_1),
	.datac(!source_packet_error_0),
	.datad(!source_ready),
	.datae(!\packet_multi:source_state.start~q ),
	.dataf(!\packet_multi:source_state.end1~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'hFFFFFDFFFFFFFFFF;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~4 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\Selector1~1_combout ),
	.datad(!\packet_multi:count_finished~combout ),
	.datae(!\source_comb_update_2~1_combout ),
	.dataf(!\Selector1~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~4 .extended_lut = "off";
defparam \Selector1~4 .lut_mask = 64'hDF8FFFFFFFFFFFFF;
defparam \Selector1~4 .shared_arith = "off";

dffeas \packet_multi:source_state.sop (
	.clk(clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_multi:source_state.sop~q ),
	.prn(vcc));
defparam \packet_multi:source_state.sop .is_wysiwyg = "true";
defparam \packet_multi:source_state.sop .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\packet_error0~combout ),
	.datac(!source_ready),
	.datad(!\packet_multi:source_state.sop~q ),
	.datae(!\packet_multi:count_finished~combout ),
	.dataf(!\packet_multi:source_state.run1~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hDFFFD5FFFFFFFFFF;
defparam \Selector2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!at_source_valid_s1),
	.datab(!\packet_error0~combout ),
	.datac(!source_ready),
	.datad(!\packet_multi:source_state.start~q ),
	.datae(!\packet_multi:source_state.end1~q ),
	.dataf(!\source_comb_update_2~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!at_source_valid_s1),
	.datab(!source_ready),
	.datac(!\Selector1~1_combout ),
	.datad(!\packet_multi:count_finished~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'hDF8FDF8FDF8FDF8F;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \at_source_valid_int~1 (
	.dataa(!at_source_valid_s1),
	.datab(!\packet_error0~combout ),
	.datac(gnd),
	.datad(!\packet_multi:count_finished~combout ),
	.datae(!\packet_multi:source_state.end1~q ),
	.dataf(!\Selector3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\at_source_valid_int~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \at_source_valid_int~1 .extended_lut = "off";
defparam \at_source_valid_int~1 .lut_mask = 64'hFFFFFFBBFFFFFFFF;
defparam \at_source_valid_int~1 .shared_arith = "off";

cyclonev_lcell_comb \at_source_valid_int~2 (
	.dataa(!at_source_valid_s1),
	.datab(!source_packet_error_1),
	.datac(!source_packet_error_0),
	.datad(!\valid_ctrl_int~q ),
	.datae(!\first_data~q ),
	.dataf(!\valid_ctrl_int1~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\at_source_valid_int~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \at_source_valid_int~2 .extended_lut = "off";
defparam \at_source_valid_int~2 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \at_source_valid_int~2 .shared_arith = "off";

cyclonev_lcell_comb \at_source_valid_int~3 (
	.dataa(!\at_source_valid_int~0_combout ),
	.datab(!\Selector2~0_combout ),
	.datac(!\Selector1~0_combout ),
	.datad(!\Selector1~2_combout ),
	.datae(!\at_source_valid_int~1_combout ),
	.dataf(!\at_source_valid_int~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\at_source_valid_int~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \at_source_valid_int~3 .extended_lut = "off";
defparam \at_source_valid_int~3 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \at_source_valid_int~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!at_source_valid_s1),
	.datab(!source_packet_error_1),
	.datac(!source_packet_error_0),
	.datad(!source_ready),
	.datae(!\packet_multi:source_state.start~q ),
	.dataf(!\packet_multi:source_state.end1~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'hFFFFFFFFFDFFFFFF;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!at_source_valid_s1),
	.datab(!\packet_error0~combout ),
	.datac(!source_ready),
	.datad(!\packet_multi:count_finished~combout ),
	.datae(!\Selector3~0_combout ),
	.dataf(!\Selector5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \Selector5~1 .shared_arith = "off";

endmodule
